** Complete Step 8: Capacitance Sweep AND Inverter Load Test
** Include model files
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45n1svt.inc'
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45p1svt.inc'
.include 'NAND_X1-post-layout.sp'

.param vdd_val=1.1
.param cap_load=5f
.TEMP 25

.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0

.vec 'input.vec'

** Power supplies
Vgnd gnd 0 0
Vsupply vdd 0 vdd_val

** Define minimum inverter subcircuit (Wn=120nm, Wp=240nm)
.subckt min_inv GND VDD IN OUT
Mp OUT IN VDD VDD g45p1svt L=45n W=240n
Mn OUT IN GND GND g45n1svt L=45n W=120n
.ends

** Main NAND gate
Xnand a b gnd vdd y NAND_X1

** Load capacitance
Cload y 0 cap_load

** PART 1: Sweep for Result 8.1 - just capacitor loads
.tran 1p 2.5n SWEEP cap_load 2f 30f 5f

** Measurements for Result 8.1
.MEASURE TRAN tpdr
+ TRIG=v(a) VAL='0.5*vdd_val' FALL=1
+ TARG=v(y) VAL='0.5*vdd_val' RISE=1

.MEASURE TRAN tpdf
+ TRIG=v(a) VAL='0.5*vdd_val' RISE=1
+ TARG=v(y) VAL='0.5*vdd_val' FALL=1

** PART 2: Add inverter load test for Result 8.2
.ALTER INVERTER_LOAD_TEST
** Set cap to 4fF
.param cap_load=4f
** No sweep this time
.tran 1p 2.5n

** Add 6 parallel minimum inverters (Wn=120nm, Wp=240nm)
** Total gate width per inverter = 360nm
Xinv1 gnd vdd y dummy1 min_inv
Xinv2 gnd vdd y dummy2 min_inv
Xinv3 gnd vdd y dummy3 min_inv
Xinv4 gnd vdd y dummy4 min_inv
Xinv5 gnd vdd y dummy5 min_inv
Xinv6 gnd vdd y dummy6 min_inv

** Measure tpdr with 4fF + 6 inverters
.MEASURE TRAN tpdr_inv_load
+ TRIG=v(a) VAL='0.5*vdd_val' FALL=1
+ TARG=v(y) VAL='0.5*vdd_val' RISE=1

.print tran v(a) v(b) v(y)
.option post
.END
