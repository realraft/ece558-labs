*
*
*
*                       LINUX           Wed Oct  1 21:15:42 2025
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 24.1.0-p089
*  Build Date     : Wed Dec 18 09:06:09 PST 2024
*
*  HSPICE LIBRARY
*
*  QRC_TECH_DIR /ece558_658/pdk/verification/qrc/typical 
*
*
*

*
.SUBCKT NAND_X1 A B GND VDD Y
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MNM0	Y#1	A#3	net13#4	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=13.0716 scb=0.0128391 scc=0.000407874 fw=2.4e-07
MNM1	net13	B#3	GND#1	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=14.2234 scb=0.0145618 scc=0.000570747 fw=2.4e-07
MPM1	Y#3	A#1	VDD#1	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=15.8854 scb=0.0156321 scc=0.000428412 fw=2.4e-07
MPM0	Y#6	B#1	VDD#3	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=17.0124 scb=0.0173035 scc=0.000589955 fw=2.4e-07
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rl1	A#1	A#2	453.826050	$poly_conn
Rl2	A#2	A#3	84.595306	$poly_conn
Rl3	B#1	B#2	351.902954	$poly_conn
Rl4	B#2	B#3	188.441467	$poly_conn
Rk1	VDD#1	VDD#2	31.000000	$metal1_conn
Rk2	Y#1	Y#2	37.500000	$metal1_conn
Rk3	A	A#2	45.164330	$metal1_conn
Rk5	Y#4	Y#7	0.410273	$metal1_conn
Rk7	Y#3	Y#4	31.000000	$metal1_conn
Rk8	Y#6	Y#7	31.000000	$metal1_conn
Rk10	net13#2	net13#5	0.408106	$metal1_conn
Rk12	net13	net13#2	37.500000	$metal1_conn
Rk13	net13#4	net13#5	37.500000	$metal1_conn
Rk14	B	B#2	45.793804	$metal1_conn
Rk15	VDD#3	VDD#4	31.000000	$metal1_conn
Rk16	GND#1	GND#2	37.500000	$metal1_conn
Rk17	Y	Y#9	0.194219	$metal1_conn
Rk18	Y#9	Y#10	0.614038	$metal1_conn
Rk19	VDD#5	VDD#7	0.107867	$metal1_conn
Rk20	VDD#7	VDD	0.059066	$metal1_conn
Rk21	VDD	VDD#8	0.044557	$metal1_conn
Rk22	VDD#6	VDD#7	18.750000	$metal1_conn
Rk23	GND#3	GND#5	0.107717	$metal1_conn
Rk24	GND#5	GND	0.055734	$metal1_conn
Rk25	GND#4	GND#5	15.500000	$metal1_conn
Rj1	VDD#8	VDD#2	0.990993	$metal2_conn
Rj2	Y#10	Y#2	1.160805	$metal2_conn
Rj3	Y#7	Y#9	1.177786	$metal2_conn
Rj4	VDD#5	VDD#4	0.988567	$metal2_conn
Rj5	GND#2	GND#3	0.990993	$metal2_conn
*
*       CAPACITOR CARDS
*
*
C1	A	B	6.9788e-18
C2	B	A#2	2.42922e-17
C3	B#1	VDD	2.7275e-17
C4	A#1	VDD	2.7618e-17
C5	Y#10	B	5.02301e-17
C6	VDD#5	VDD	5.6948e-17
C7	VDD#4	VDD	1.6529e-17
C8	A#1	B#1	4.44092e-18
C9	Y	VDD#4	4.27623e-18
C10	Y#9	VDD	2.60906e-18
C11	VDD#8	VDD	5.06912e-17
C12	A#1	B#2	1.05094e-18
C13	A#3	B#3	1.81005e-18
C14	VDD#5	B#1	4.84004e-18
C15	VDD#2	VDD	1.54934e-17
C16	VDD#4	B#1	6.17036e-18
C17	A#2	B#3	1.99786e-18
C18	VDD#4	A#1	5.79241e-19
C19	Y#9	B#1	9.07265e-19
C20	VDD#6	VDD	2.51287e-17
C21	A#2	B#2	6.09814e-18
C22	GND#2	B#3	6.17036e-18
C23	Y#9	A#1	1.28235e-18
C24	GND#3	B#3	4.23041e-18
C25	VDD#2	B#1	6.23537e-19
C26	GND#3	B#2	2.03135e-18
C27	VDD#8	A#1	4.97748e-18
C28	VDD#4	VDD#5	8.62319e-18
C29	VDD#2	A#1	6.16783e-18
C30	Y#9	B#2	7.94046e-17
C31	Y#9	A#2	1.23595e-18
C32	Y#2	B#3	6.03619e-19
C33	VDD#6	B#1	8.90318e-19
C34	GND#3	GND#2	8.03771e-18
C35	Y#2	A#3	6.07448e-18
C36	GND#4	B#3	6.88567e-19
C37	B#2	Y#10	5.3079e-18
C38	VDD#6	A#1	7.57109e-19
C39	Y#10	A#2	1.94415e-17
C40	Y#2	A#2	1.6535e-17
C41	VDD#4	VDD#3	4.92159e-18
C42	GND#2	GND#4	2.291e-18
C43	VDD#5	VDD#6	5.719e-19
C44	Y#10	Y#9	3.7233e-18
C45	GND#3	GND#4	8.80726e-19
C46	VDD#4	VDD#6	2.37993e-18
C47	GND#2	GND#1	4.92159e-18
C48	VDD#2	VDD#8	8.41881e-18
C49	Y#10	VDD#2	4.09523e-18
C50	VDD#2	VDD#1	4.92159e-18
C51	VDD#8	VDD#6	5.85256e-19
C52	VDD#2	VDD#6	2.46733e-18
C53	Y#2	Y#1	4.92159e-18
C54	Y#4	Y#3	2.07801e-18
C55	GND#3	GND	5.8791e-17
C56	Y#9	Y#7	4.80932e-18
C57	Y#4	A#1	4.32919e-18
C58	net13#5	B#3	6.65212e-19
C59	Y#4	Y#7	1.18344e-17
C60	GND#3	net13#2	1.24427e-17
C61	Y#7	VDD#5	1.22482e-17
C62	net13#2	B#2	1.06392e-17
C63	Y#10	Y#4	6.37156e-18
C64	Y#7	A#1	2.51541e-18
C65	Y#4	VDD#6	1.31981e-17
C66	net13#5	Y#10	7.9664e-19
C67	Y#7	Y#6	2.20949e-18
C68	GND#4	net13#2	1.33315e-17
C69	net13#5	B#2	2.89881e-18
C70	net13#2	Y#9	2.56364e-18
C71	net13#5	net13#4	1.96797e-18
C72	net13#5	net13#2	8.76265e-18
C73	Y#4	B#1	7.8168e-19
C74	net13#2	GND#2	5.28939e-17
C75	VDD#2	Y#4	5.28731e-17
C76	Y#7	B#1	6.92763e-18
C77	net13#2	net13	1.95976e-18
C78	Y#4	B	6.46005e-19
C79	Y#7	VDD#4	5.64394e-17
C80	GND#4	GND	2.54356e-17
C81	GND#4	net13#5	1.26489e-17
C82	Y#9	Y#4	1.48819e-18
C83	Y#7	VDD#6	1.57835e-17
C84	Y#4	VDD	2.68381e-17
C85	net13#5	B	7.65471e-18
C86	Y#2	net13#5	5.28731e-17
C87	Y#7	VDD	1.98157e-17
C88	GND#2	GND	1.70825e-17
C89	VDD#2	Y#7	9.64389e-19
C90	net13#2	B#3	4.33329e-18
C91	A	GND	1.29818e-17
C92	B	GND	1.9933e-17
C93	Y	GND	1.94219e-17
C94	B#1	GND	1.11619e-18
C95	A#1	GND	8.24277e-18
C96	B#3	GND	2.01593e-17
C97	A#3	GND	2.27223e-17
C98	B#2	GND	6.81979e-17
C99	A#2	GND	4.31399e-17
C100	VDD#5	GND	2.48168e-19
C101	VDD#4	GND	5.37996e-19
C102	Y#9	GND	2.39668e-17
C103	Y#10	GND	2.65796e-17
C104	Y#2	GND	3.10959e-17
C105	net13#2	GND	1.04592e-17
C106	net13#5	GND	2.89669e-17
*
*
.ENDS NAND_X1
*
