*
*
*
*                       LINUX           Sun Oct 19 14:43:58 2025
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 24.1.0-p089
*  Build Date     : Wed Dec 18 09:06:09 PST 2024
*
*  HSPICE LIBRARY
*
*  QRC_TECH_DIR /ece558_658/pdk/verification/qrc/typical 
*
*
*

*
.SUBCKT HA_ACCUM A! B! CIN COUT GND PHI PHI! RST SOUT VDD
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MXI0/XI0/XI0/MNM0	A!#7	CIN#3	GND#1	GND	g45n1svt
+ L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.90867 scb=0.00164474 scc=3.75172e-06 fw=1.2e-07
MXI1/XI5/MNM0	XI1/D#5	RST#1	XI1/XI5/net13#4	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.82604 scb=0.000193838 scc=1.85478e-08 fw=2.4e-07
MXI1/XI4/XI1/MNM0	PHI!#7	PHI#3	GND#3	GND	g45n1svt
+ L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.99885 scb=0.00021225 scc=1.92763e-08 fw=1.2e-07
MXI0/XI0/XI1/MNM0	B!#8	SOUT#3	GND#5	GND	g45n1svt
+ L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI1/XI5/MNM1	XI1/XI5/net13	net3	GND#7	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI1/XI0/MNM1	XI0/XI1/XI0/net13#5	SOUT#4	GND#9	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI4/MNM0	XI1/XI4/net24#5	PHI!#3	XI1/XI4/net36	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI4/MNM3	XI1/XI4/net36	XI1/D	GND#11	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI0/MNM2	XI0/XI0/net15	B!#1	GND#13	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI0/XI0/MNM0	net3#17	A!#3	XI0/XI0/net15	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI0/XI1/XI0/MNM0	XI0/XI1/net2#10	CIN#4	XI0/XI1/XI0/net13
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI4/MNM2	XI1/XI4/net25	XI1/XI4/net24#3	GND#15	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI4/MNM1	XI1/Q#8	PHI#6	XI1/XI4/net25	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI0/MNM1	net3#13	CIN#9	XI0/XI0/net18	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI1/XI6/MNM0	SOUT#17	XI1/Q#3	GND#17	GND	g45n1svt
+ L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI0/XI0/MNM3	XI0/XI0/net18	SOUT#9	GND#21	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI0/XI1/XI2/MNM0	COUT#4	XI0/XI1/net2	GND#19	GND	g45n1svt
+ L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI0/XI0/XI0/MPM0	A!#5	CIN#1	VDD#1	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.95118 scb=0.00508612 scc=7.502e-05 fw=2.4e-07
MXI1/XI5/MPM1	XI1/D#11	RST#3	VDD#6	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.26407 scb=0.00404065 scc=4.42753e-05 fw=2.4e-07
MXI1/XI4/XI1/MPM0	PHI!#5	PHI#1	VDD#3	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.1139 scb=0.00244911 scc=5.96896e-06 fw=2.4e-07
MXI0/XI0/XI1/MPM0	B!#6	SOUT#1	VDD#7	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI1/XI5/MPM0	XI1/D#8	net3#3	VDD#9	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI0/XI1/XI0/MPM0	XI0/XI1/net2#7	SOUT#6	VDD#11	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI1/XI4/MPM3	XI1/Q#4	PHI!#1	XI1/XI4/net17	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI1/XI4/MPM2	XI1/XI4/net17	XI1/XI4/net24	VDD#13	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI0/XI0/MPM0	XI0/XI0/net4	SOUT#7	VDD#15	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI0/XI0/MPM1	net3#10	A!#1	XI0/XI0/net4	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI0/XI1/XI0/MPM1	XI0/XI1/net2#4	CIN#6	VDD#19	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI1/XI4/MPM0	XI1/XI4/net9	XI1/D#3	VDD#17	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI1/XI4/MPM1	XI1/XI4/net24#10	PHI#4	XI1/XI4/net9	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI0/XI0/MPM3	net3#7	CIN#7	XI0/XI0/net11	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI1/XI6/MPM0	SOUT#15	XI1/Q	VDD#21	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
MXI0/XI0/MPM2	XI0/XI0/net11	B!#3	VDD#25	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI0/XI1/XI2/MPM0	COUT#2	XI0/XI1/net2#3	VDD#23	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 fw=2.4e-07
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rl1	CIN#1	CIN#2	306.867249	$poly_conn
Rl2	CIN#2	CIN#3	383.790314	$poly_conn
Rl3	RST#1	RST#2	76.098015	$poly_conn
Rl4	RST#2	RST#3	606.867249	$poly_conn
Rl5	PHI#1	PHI#2	199.979935	$poly_conn
Rl6	PHI#2	PHI#3	492.287628	$poly_conn
Rl7	SOUT#1	SOUT#2	142.287613	$poly_conn
Rl8	SOUT#2	SOUT#3	549.979919	$poly_conn
Rl9	net3	net3#2	622.251892	$poly_conn
Rl10	net3#2	net3#3	60.713398	$poly_conn
Rl11	SOUT#4	SOUT#5	215.364548	$poly_conn
Rl12	SOUT#5	SOUT#6	469.210693	$poly_conn
Rl13	PHI!#1	PHI!#2	206.461472	$poly_conn
Rl14	PHI!#2	PHI!#3	391.076874	$poly_conn
Rl15	XI1/XI4/net24	XI1/XI4/net24#2	490.321899	$poly_conn
Rl16	XI1/D	XI1/D#2	117.244949	$poly_conn
Rl17	SOUT#7	SOUT#8	101.860336	$poly_conn
Rl18	B!#1	B!#2	141.475723	$poly_conn
Rl19	A!#1	A!#2	372.251862	$poly_conn
Rl20	A!#2	A!#3	210.713394	$poly_conn
Rl21	CIN#4	CIN#5	418.405701	$poly_conn
Rl22	CIN#5	CIN#6	264.559540	$poly_conn
Rl23	XI1/D#3	XI1/D#4	53.014187	$poly_conn
Rl24	XI1/XI4/net24#3	XI1/XI4/net24#4	145.321869
+ $poly_conn
Rl25	PHI#4	PHI#5	126.098015	$poly_conn
Rl26	PHI#5	PHI#6	464.559570	$poly_conn
Rl27	CIN#7	CIN#8	222.251862	$poly_conn
Rl28	CIN#8	CIN#9	360.713379	$poly_conn
Rl29	XI1/Q	XI1/Q#2	449.174927	$poly_conn
Rl30	XI1/Q#2	XI1/Q#3	241.482620	$poly_conn
Rl31	XI0/XI1/net2	XI0/XI1/net2#2	560.713379	$poly_conn
Rl32	XI0/XI1/net2#2	XI0/XI1/net2#3	129.944168	$poly_conn
Rl33	B!#3	B!#4	60.706493	$poly_conn
Rl34	SOUT#9	SOUT#10	113.398796	$poly_conn
Rk1	VDD#1	VDD#2	31.000000	$metal1_conn
Rk2	GND#1	GND#2	75.000000	$metal1_conn
Rk3	XI1/D#5	XI1/D#6	37.501156	$metal1_conn
Rk4	VDD#3	VDD#4	31.000000	$metal1_conn
Rk5	VDD#5	VDD#6	31.001158	$metal1_conn
Rk6	GND#3	GND#4	75.000000	$metal1_conn
Rk7	A!#4	A!#5	31.001158	$metal1_conn
Rk8	A!#6	A!#7	75.001549	$metal1_conn
Rk9	PHI!#4	PHI!#5	31.001158	$metal1_conn
Rk10	PHI!#6	PHI!#7	75.001549	$metal1_conn
Rk11	VDD#7	VDD#8	31.000000	$metal1_conn
Rk12	XI1/XI5/net13#2	XI1/XI5/net13#3	0.001157
+ $metal1_conn
Rk13	XI1/XI5/net13#3	XI1/XI5/net13#5	0.232308
+ $metal1_conn
Rk15	XI1/XI5/net13	XI1/XI5/net13#2	37.500000	$metal1_conn
Rk16	XI1/XI5/net13#4	XI1/XI5/net13#5	37.500000
+ $metal1_conn
Rk17	GND#5	GND#6	75.000000	$metal1_conn
Rk18	XI1/D#7	XI1/D#9	0.001157	$metal1_conn
Rk19	XI1/D#9	XI1/D#10	0.120231	$metal1_conn
Rk20	XI1/D#10	XI1/D#12	0.114924	$metal1_conn
Rk22	XI1/D#8	XI1/D#9	31.000000	$metal1_conn
Rk23	XI1/D#11	XI1/D#12	31.000000	$metal1_conn
Rk24	B!#5	B!#6	31.001158	$metal1_conn
Rk25	GND#7	GND#8	37.500000	$metal1_conn
Rk26	VDD#9	VDD#10	31.000000	$metal1_conn
Rk27	B!#7	B!#8	75.001549	$metal1_conn
Rk28	XI1/D#14	XI1/D#15	0.450092	$metal1_conn
Rk29	XI1/D#15	XI1/D#16	0.266916	$metal1_conn
Rk30	GND#9	GND#10	37.500000	$metal1_conn
Rk31	VDD#11	VDD#12	31.000000	$metal1_conn
Rk32	XI1/Q#4	XI1/Q#5	15.500000	$metal1_conn
Rk33	XI1/XI4/net24#5	XI1/XI4/net24#6	37.500000
+ $metal1_conn
Rk34	PHI!#2	PHI!	45.682796	$metal1_conn
Rk35	PHI!	PHI!#9	0.833515	$metal1_conn
Rk36	VDD#13	VDD#14	15.500000	$metal1_conn
Rk37	GND#11	GND#12	37.500000	$metal1_conn
Rk38	VDD#15	VDD#16	15.500000	$metal1_conn
Rk39	GND#13	GND#14	37.500000	$metal1_conn
Rk40	XI1/Q#6	XI1/Q#7	0.365328	$metal1_conn
Rk41	A!#2	A!	45.478970	$metal1_conn
Rk42	A!	A!#9	1.376578	$metal1_conn
Rk44	XI0/XI1/XI0/net13#2	XI0/XI1/XI0/net13#4	0.232308
+ $metal1_conn
Rk45	XI0/XI1/XI0/net13#4	XI0/XI1/XI0/net13#5	37.501156
+ $metal1_conn
Rk46	XI0/XI1/XI0/net13	XI0/XI1/XI0/net13#2	37.500000
+ $metal1_conn
Rk48	XI0/XI1/net2#5	XI0/XI1/net2#8	0.237615	$metal1_conn
Rk49	XI0/XI1/net2#8	XI0/XI1/net2#9	0.001157	$metal1_conn
Rk50	XI0/XI1/net2#4	XI0/XI1/net2#5	31.000000	$metal1_conn
Rk51	XI0/XI1/net2#7	XI0/XI1/net2#8	31.000000	$metal1_conn
Rk52	XI1/D#17	XI1/D#2	0.292025	$metal1_conn
Rk53	XI1/D#2	XI1/D#19	0.466581	$metal1_conn
Rk54	CIN#5	CIN#11	45.731133	$metal1_conn
Rk55	SOUT#11	SOUT#8	0.156463	$metal1_conn
Rk56	SOUT#8	SOUT#2	45.836899	$metal1_conn
Rk57	VDD#17	VDD#18	15.500000	$metal1_conn
Rk58	GND#15	GND#16	37.500000	$metal1_conn
Rk59	VDD#19	VDD#20	31.001158	$metal1_conn
Rk60	XI1/XI4/net24#4	XI1/XI4/net24#2	45.402275
+ $metal1_conn
Rk61	XI1/XI4/net24#2	XI1/XI4/net24#9	0.668824
+ $metal1_conn
Rk62	XI1/D#20	XI1/D#4	45.082287	$metal1_conn
Rk63	XI1/XI4/net24#10	XI1/XI4/net24#11	15.500000
+ $metal1_conn
Rk64	XI1/XI4/net24#12	XI1/XI4/net24#13	0.688239
+ $metal1_conn
Rk65	XI1/Q#8	XI1/Q#9	37.500000	$metal1_conn
Rk66	XI0/XI1/net2#11	XI0/XI1/net2#12	0.001157
+ $metal1_conn
Rk67	XI0/XI1/net2#12	XI0/XI1/net2#13	0.169876
+ $metal1_conn
Rk68	XI0/XI1/net2#10	XI0/XI1/net2#11	37.500000
+ $metal1_conn
Rk69	net3#4	net3#2	46.295746	$metal1_conn
Rk70	B!#9	B!	1.630869	$metal1_conn
Rk71	B!	B!#10	1.130727	$metal1_conn
Rk72	B!#11	B!#2	45.782852	$metal1_conn
Rk74	net3#6	net3#9	0.322022	$metal1_conn
Rk75	net3#9	net3#11	0.257371	$metal1_conn
Rk77	net3#7	net3#6	15.500000	$metal1_conn
Rk78	net3#10	net3#11	15.500000	$metal1_conn
Rk80	net3#14	net3#16	0.305642	$metal1_conn
Rk81	net3#16	net3#18	0.240992	$metal1_conn
Rk83	net3#13	net3#14	37.500000	$metal1_conn
Rk84	net3#17	net3#18	37.500000	$metal1_conn
Rk85	CIN	CIN#12	0.415576	$metal1_conn
Rk86	CIN#12	CIN#13	0.688033	$metal1_conn
Rk87	CIN#13	CIN#8	46.508373	$metal1_conn
Rk88	VDD#21	VDD#22	31.000000	$metal1_conn
Rk89	VDD#23	VDD#24	31.000000	$metal1_conn
Rk90	GND#17	GND#18	75.000000	$metal1_conn
Rk91	GND#19	GND#20	75.000000	$metal1_conn
Rk92	XI1/Q#2	XI1/Q#11	45.453136	$metal1_conn
Rk93	XI1/Q#11	XI1/Q#12	0.376483	$metal1_conn
Rk94	XI0/XI1/net2#2	XI0/XI1/net2#15	45.440205	$metal1_conn
Rk95	XI0/XI1/net2#15	XI0/XI1/net2#16	0.343778
+ $metal1_conn
Rk96	B!#4	B!#14	45.156464	$metal1_conn
Rk97	SOUT#14	SOUT#15	31.001158	$metal1_conn
Rk98	VDD#25	VDD#26	15.500000	$metal1_conn
Rk99	GND#21	GND#22	37.500000	$metal1_conn
Rk100	COUT#1	COUT#2	31.001158	$metal1_conn
Rk101	SOUT#16	SOUT#17	75.001549	$metal1_conn
Rk102	COUT#3	COUT#4	75.001549	$metal1_conn
Rk103	SOUT#18	SOUT#19	1.205139	$metal1_conn
Rk104	SOUT#20	SOUT#5	46.880508	$metal1_conn
Rk105	SOUT#22	SOUT#10	0.248977	$metal1_conn
Rk106	SOUT#10	SOUT#24	0.776813	$metal1_conn
Rk107	COUT#5	COUT#6	0.885980	$metal1_conn
Rk108	VDD#27	VDD#29	0.045855	$metal1_conn
Rk109	VDD#29	VDD#30	0.256720	$metal1_conn
Rk110	VDD#30	VDD#31	0.194163	$metal1_conn
Rk111	VDD#31	VDD#32	0.085599	$metal1_conn
Rk112	VDD#32	VDD#33	0.390413	$metal1_conn
Rk113	VDD#33	VDD	0.104388	$metal1_conn
Rk114	VDD#28	VDD#29	18.750000	$metal1_conn
Rk115	VDD#34	VDD#36	0.047483	$metal1_conn
Rk116	VDD#36	VDD#37	0.214504	$metal1_conn
Rk117	VDD#37	VDD#38	0.041755	$metal1_conn
Rk118	VDD#38	VDD#39	0.185811	$metal1_conn
Rk119	VDD#39	VDD#40	0.085599	$metal1_conn
Rk120	VDD#40	VDD#41	0.081423	$metal1_conn
Rk121	VDD#41	VDD#42	0.151363	$metal1_conn
Rk122	VDD#42	VDD#43	0.044887	$metal1_conn
Rk123	VDD#43	VDD#44	0.125266	$metal1_conn
Rk124	VDD#44	VDD	0.114827	$metal1_conn
Rk125	VDD#35	VDD#36	18.750000	$metal1_conn
Rk126	GND#23	GND#25	0.156403	$metal1_conn
Rk127	GND#25	GND#26	0.045855	$metal1_conn
Rk128	GND#26	GND#27	0.167022	$metal1_conn
Rk129	GND#27	GND#28	0.313165	$metal1_conn
Rk130	GND#28	GND#29	0.277673	$metal1_conn
Rk131	GND#29	GND#30	0.129442	$metal1_conn
Rk132	GND#30	GND	0.119003	$metal1_conn
Rk133	GND#24	GND#25	15.500000	$metal1_conn
Rk134	COUT	COUT#7	0.671134	$metal1_conn
Rk135	PHI#7	PHI#8	1.759981	$metal1_conn
Rk136	PHI#8	PHI#9	1.695851	$metal1_conn
Rk137	PHI#9	PHI	0.454367	$metal1_conn
Rk138	RST#4	RST#5	3.362283	$metal1_conn
Rk139	RST#5	RST	0.414858	$metal1_conn
Rk140	GND#31	GND#32	15.548018	$metal1_conn
Rk141	GND#32	GND#33	0.210865	$metal1_conn
Rk142	GND#33	GND#34	0.194163	$metal1_conn
Rk143	GND#34	GND#35	0.085599	$metal1_conn
Rk144	GND#35	GND#36	0.070984	$metal1_conn
Rk145	GND#36	GND#37	0.151363	$metal1_conn
Rk146	GND#37	GND#38	0.168065	$metal1_conn
Rk147	GND#38	GND	0.104388	$metal1_conn
Rk166	PHI#5	PHI#8	45.000000	$metal1_conn
Rk167	PHI#2	PHI#9	45.000000	$metal1_conn
Rk168	RST#2	RST#5	45.000000	$metal1_conn
Rk159	CIN#2	CIN#12	45.000000	$metal1_conn
Rj1	GND#2	GND#30	1.223605	$metal2_conn
Rj2	XI1/D#6	XI1/D#16	1.048436	$metal2_conn
Rj3	VDD#33	VDD#4	0.993049	$metal2_conn
Rj4	GND#4	GND#38	1.209022	$metal2_conn
Rj5	VDD#2	VDD#48	0.480633	$metal2_conn
Rj6	VDD#48	VDD#5	0.464040	$metal2_conn
Rj7	A!#4	A!#9	0.906232	$metal2_conn
Rj8	A!#9	A!#6	0.845129	$metal2_conn
Rj9	PHI!#4	PHI!#9	0.677766	$metal2_conn
Rj10	PHI!#9	PHI!#6	1.073595	$metal2_conn
Rj11	XI1/D#15	XI1/D#10	1.727739	$metal2_conn
Rj12	VDD#43	VDD#8	0.983327	$metal2_conn
Rj13	GND#6	GND#29	1.223605	$metal2_conn
Rj14	B!#5	B!#10	0.813873	$metal2_conn
Rj15	B!#10	B!#7	0.937488	$metal2_conn
Rj16	GND#37	GND#8	0.968744	$metal2_conn
Rj17	VDD#10	VDD#42	0.970427	$metal2_conn
Rj18	XI1/D#19	XI1/D#14	1.904141	$metal2_conn
Rj19	CIN#11	CIN#13	2.331907	$metal2_conn
Rj20	GND#36	GND#10	0.968744	$metal2_conn
Rj21	VDD#12	VDD#41	0.970427	$metal2_conn
Rj22	XI1/Q#5	XI1/Q#7	0.829161	$metal2_conn
Rj23	XI1/XI4/net24#13	XI1/XI4/net24#9	0.692283
+ $metal2_conn
Rj24	XI1/XI4/net24#9	XI1/XI4/net24#6	0.510336
+ $metal2_conn
Rj25	VDD#32	VDD#14	0.902076	$metal2_conn
Rj26	GND#12	GND#35	0.968744	$metal2_conn
Rj27	VDD#40	VDD#16	0.906937	$metal2_conn
Rj28	GND#14	GND#28	0.973605	$metal2_conn
Rj29	XI1/Q#6	XI1/Q#12	1.453691	$metal2_conn
Rj30	XI0/XI1/net2#16	XI0/XI1/net2#5	1.014175	$metal2_conn
Rj31	XI1/D#20	XI1/D#17	1.637058	$metal2_conn
Rj32	SOUT#11	SOUT#24	1.578456	$metal2_conn
Rj33	VDD#31	VDD#18	0.902076	$metal2_conn
Rj34	GND#16	GND#34	0.968744	$metal2_conn
Rj35	VDD#20	VDD#39	0.970427	$metal2_conn
Rj36	XI1/XI4/net24#11	XI1/XI4/net24#12	1.125680
+ $metal2_conn
Rj37	XI1/Q#11	XI1/Q#9	1.099990	$metal2_conn
Rj38	XI0/XI1/net2#13	XI0/XI1/net2#15	1.758312
+ $metal2_conn
Rj39	net3#4	net3#23	1.156232	$metal2_conn
Rj40	net3#23	net3#16	1.452751	$metal2_conn
Rj41	B!#14	B!#9	0.801380	$metal2_conn
Rj42	B!#9	B!#11	0.679856	$metal2_conn
Rj43	VDD#30	VDD#22	0.993049	$metal2_conn
Rj44	GND#20	GND#56	0.726111	$metal2_conn
Rj45	GND#56	GND#18	0.704161	$metal2_conn
Rj46	VDD#24	VDD#38	0.988998	$metal2_conn
Rj47	SOUT#14	SOUT#19	1.115254	$metal2_conn
Rj48	SOUT#19	SOUT#16	0.636107	$metal2_conn
Rj49	VDD#37	VDD#26	0.907747	$metal2_conn
Rj50	GND#22	GND#27	0.973605	$metal2_conn
Rj51	COUT#3	COUT#6	0.757632	$metal2_conn
Rj52	COUT#6	COUT#1	0.993729	$metal2_conn
Rj53	SOUT	SOUT#18	1.273576	$metal2_conn
Rj54	SOUT#18	SOUT#20	0.921903	$metal2_conn
Rj55	SOUT#20	SOUT#22	2.500540	$metal2_conn
Rj56	COUT#5	COUT#7	2.725023	$metal2_conn
Rj57	GND#32	GND#26	3.882558	$metal2_conn
Rj58	VDD#27	VDD#34	3.921446	$metal2_conn
Rj141	net3#9	net3#23	0.500000	$metal2_conn
Rj151	GND#33	GND#56	0.500000	$metal2_conn
Rj68	VDD#44	VDD#48	0.500000	$metal2_conn
*
*       CAPACITOR CARDS
*
*
C1	VDD#39	CIN#6	4.16751e-18
C2	net3#16	A!#2	2.38906e-18
C3	COUT#6	SOUT#20	8.74186e-17
C4	XI1/XI4/net24#4	XI1/Q#11	1.49839e-17
C5	VDD#20	CIN#6	4.0872e-18
C6	VDD#16	net3#9	2.69354e-18
C7	VDD#34	GND#31	1.39542e-17
C8	COUT#6	XI0/XI1/net2	7.48119e-18
C9	SOUT#18	XI1/Q#3	1.55626e-18
C10	CIN#11	SOUT#5	2.7909e-17
C11	VDD#18	XI1/D#3	6.45552e-18
C12	SOUT#10	CIN#8	3.40191e-18
C13	PHI!#6	XI1/D#19	8.36117e-18
C14	XI1/XI4/net24#6	XI1/D	1.8988e-18
C15	VDD#44	RST#3	4.10956e-18
C16	COUT#3	XI0/XI1/net2	5.18165e-18
C17	VDD#31	XI1/D#3	4.10481e-18
C18	RST#2	CIN#4	1.53357e-17
C19	COUT#3	SOUT#20	1.99738e-17
C20	XI1/D#2	PHI!#3	3.94365e-17
C21	XI1/XI4/net24#12	XI1/XI4/net24#4	1.1037e-18
C22	XI1/D#19	XI1/XI4/net24#9	4.53836e-18
C23	VDD#41	net3#2	9.35443e-18
C24	CIN#8	B!#4	3.19507e-18
C25	XI1/D#14	SOUT#5	7.88532e-18
C26	GND#34	GND#16	1.0238e-17
C27	VDD#43	VDD#42	1.68608e-17
C28	B!#5	B!#6	8.47836e-18
C29	net3#9	A!#1	1.29015e-18
C30	VDD#40	net3#9	1.69894e-18
C31	XI1/XI4/net24#2	PHI!#3	1.97764e-17
C32	XI1/D#17	XI1/Q#9	7.80585e-18
C33	SOUT#20	XI0/XI1/net2	2.18236e-17
C34	GND#28	GND#14	9.66245e-18
C35	VDD#18	PHI#4	2.37746e-18
C36	XI1/D#10	CIN#11	1.24968e-17
C37	B!#2	B!#9	8.98145e-18
C38	VDD#12	net3#2	1.29263e-17
C39	VDD#31	PHI#4	4.96959e-18
C40	VDD#27	GND#31	1.79196e-17
C41	XI1/Q#5	XI1/Q#4	9.30041e-18
C42	net3#4	CIN#5	1.24619e-17
C43	XI1/D#19	XI1/XI4/net24#6	1.52085e-17
C44	XI1/Q#11	PHI#5	1.16343e-17
C45	XI1/XI4/net24#11	XI1/XI4/net24#10	7.53548e-18
C46	XI1/XI4/net24#11	XI1/D#4	3.45102e-18
C47	SOUT#5	CIN#4	4.20801e-18
C48	net3#4	CIN#6	1.35025e-17
C49	GND#12	PHI!#3	2.02958e-18
C50	XI1/D#17	XI1/Q#11	1.88368e-17
C51	SOUT#10	B!#4	2.61929e-18
C52	XI1/XI4/net24#11	XI1/D#3	3.27281e-18
C53	VDD#27	XI1/Q#3	1.24354e-18
C54	A!#4	CIN#1	6.05749e-18
C55	XI0/XI1/net2#15	CIN#5	7.43893e-18
C56	XI1/XI4/net24#12	PHI#5	4.06087e-17
C57	net3#9	VDD#38	7.00273e-18
C58	XI1/D#15	CIN#11	5.94265e-18
C59	SOUT#22	COUT#7	1.19535e-16
C60	XI1/D#19	PHI!#2	5.57418e-18
C61	VDD#5	RST#3	5.42714e-18
C62	GND#32	XI0/XI1/net2	1.0422e-18
C63	VDD#27	PHI#7	2.49545e-17
C64	GND#35	XI1/D	2.42413e-18
C65	XI1/XI4/net24#11	PHI#5	1.50188e-17
C66	GND#10	GND#36	1.0238e-17
C67	GND#4	GND#3	3.1639e-18
C68	B!#2	A!#3	9.13179e-18
C69	XI1/XI4/net24#11	PHI#4	7.57347e-18
C70	VDD#34	XI0/XI1/net2	8.86371e-19
C71	XI1/D#17	XI1/XI4/net24#12	8.06775e-18
C72	net3#4	VDD#38	1.36924e-18
C73	SOUT#20	COUT#7	2.64737e-17
C74	GND#12	XI1/D	3.7665e-18
C75	XI1/D#2	XI1/XI4/net24#3	1.40726e-18
C76	COUT#7	VDD#35	7.44569e-18
C77	XI1/Q#6	VDD#14	1.63056e-17
C78	VDD#4	PHI#1	6.76392e-18
C79	XI1/Q#11	XI1/Q#2	3.35663e-18
C80	XI1/D#19	XI1/D#2	1.57987e-18
C81	VDD#33	PHI#1	4.6061e-18
C82	XI1/D#15	XI1/D#14	4.55699e-18
C83	GND#30	CIN#3	3.66677e-18
C84	B!#10	A!#2	1.45297e-18
C85	SOUT#20	COUT#5	1.77608e-16
C86	SOUT#22	GND#26	2.22433e-17
C87	GND#32	COUT#3	1.33266e-18
C88	VDD#38	XI0/XI1/net2#15	3.53013e-18
C89	net3#4	VDD#24	8.36933e-18
C90	XI1/D#20	XI1/XI4/net24#12	1.96826e-17
C91	XI1/XI4/net24#12	XI1/Q#2	2.89847e-18
C92	GND#2	CIN#3	3.96405e-18
C93	GND#27	net3#16	9.27251e-18
C94	XI1/D#6	GND#38	1.65558e-17
C95	A!#6	GND#6	1.4863e-17
C96	XI1/Q#6	VDD#32	4.14214e-18
C97	GND#30	A!#6	1.31853e-17
C98	VDD#18	VDD#31	1.16687e-17
C99	net3#9	CIN#8	1.55592e-17
C100	CIN#13	VDD#8	6.29073e-18
C101	XI1/XI4/net24#11	XI1/Q	4.03173e-18
C102	CIN#3	SOUT#3	7.17245e-18
C103	XI1/Q#9	SOUT#16	1.50349e-18
C104	CIN#2	VDD#2	3.99391e-18
C105	XI1/D#20	XI1/XI4/net24#11	1.3057e-17
C106	SOUT#20	GND#32	1.25561e-17
C107	CIN#1	SOUT#2	2.69766e-18
C108	XI1/XI4/net24#9	PHI!#2	1.74823e-18
C109	VDD#16	VDD#40	1.0979e-17
C110	XI0/XI1/net2#16	net3#4	3.40342e-17
C111	VDD#10	VDD#9	7.83801e-18
C112	VDD#8	CIN#1	1.73636e-18
C113	GND#28	B!#1	2.7139e-18
C114	XI1/D#10	RST#3	3.88703e-18
C115	GND#6	A!#9	5.65589e-18
C116	VDD#20	XI0/XI1/net2#3	1.01229e-18
C117	RST#1	net3	3.14306e-18
C118	CIN#13	SOUT#8	2.94542e-17
C119	GND#35	XI1/D#17	1.58396e-18
C120	B!#14	CIN#7	1.32694e-17
C121	XI1/Q#9	SOUT#19	5.36449e-18
C122	GND#26	COUT#7	1.03032e-16
C123	XI1/D#15	RST#3	1.25112e-18
C124	SOUT#18	GND#32	3.44046e-17
C125	GND#14	B!#1	4.9463e-18
C126	GND#2	A!#6	4.04959e-17
C127	GND#36	XI1/D#2	3.24657e-18
C128	VDD#43	CIN#13	3.05188e-18
C129	XI1/XI4/net24#4	PHI#6	3.61375e-17
C130	PHI#7	VDD	4.1237e-17
C131	VDD#2	VDD#1	4.59183e-18
C132	RST#3	net3#2	1.10422e-17
C133	A!#4	SOUT#1	1.96312e-18
C134	GND#36	XI1/XI4/net24#6	1.96676e-17
C135	XI0/XI1/net2#13	GND#20	1.11215e-17
C136	COUT#7	GND#32	1.43822e-17
C137	XI0/XI1/net2#16	XI0/XI1/net2#15	7.04611e-18
C138	GND#6	GND#5	3.06513e-18
C139	VDD#26	VDD#25	1.35961e-17
C140	XI1/XI4/net24#13	PHI!#2	2.64065e-17
C141	XI1/Q#11	SOUT#19	7.01749e-18
C142	PHI!#4	PHI#1	8.09825e-18
C143	XI1/XI4/net24#9	XI1/D#2	3.0624e-17
C144	GND#28	A!#3	4.34667e-18
C145	RST#4	GND#33	1.51603e-17
C146	GND#34	XI1/Q#9	1.24572e-17
C147	B!#11	CIN#8	1.64202e-18
C148	net3#9	VDD#26	2.27362e-18
C149	net3#16	SOUT#10	4.33498e-18
C150	GND#26	VDD#35	1.53511e-17
C151	net3#4	XI0/XI1/net2#2	9.28475e-19
C152	GND#33	GND#18	9.30871e-18
C153	GND#14	A!#3	2.55369e-18
C154	CIN#13	A!#2	1.52499e-17
C155	GND#20	GND#19	3.25792e-18
C156	XI1/D#17	PHI!#3	8.962e-19
C157	B!#5	VDD#42	1.54612e-17
C158	XI1/Q#7	PHI!#2	9.18965e-19
C159	COUT#5	GND#32	1.08101e-16
C160	XI1/XI4/net24#6	XI1/D#2	9.87705e-18
C161	GND#38	GND#4	9.24934e-18
C162	SOUT#18	VDD#27	2.23434e-17
C163	B!#9	CIN#8	8.66258e-17
C164	XI1/XI4/net24#12	SOUT#19	5.53384e-18
C165	VDD#44	VDD#5	1.02424e-17
C166	net3#4	XI0/XI1/net2#3	1.41355e-18
C167	VDD#38	CIN#7	3.76854e-18
C168	XI0/XI1/net2#15	XI0/XI1/net2#2	6.41939e-18
C169	PHI#6	XI1/Q#2	2.86362e-18
C170	XI1/D#6	RST#1	5.54809e-18
C171	GND#16	XI1/Q#9	3.29714e-17
C172	XI1/D#16	RST#2	5.30268e-17
C173	net3#9	VDD#37	1.33783e-18
C174	CIN#8	B!#14	8.83203e-18
C175	VDD#22	XI1/Q	4.68876e-18
C176	XI1/XI4/net24#9	XI1/XI4/net24#2	7.14446e-18
C177	VDD#34	COUT#5	1.42169e-18
C178	SOUT#8	VDD#41	7.25049e-18
C179	VDD#30	XI1/Q	4.97335e-18
C180	GND#38	RST#1	2.53688e-18
C181	XI1/XI4/net24#12	SOUT#14	3.0753e-18
C182	RST#2	XI1/D#6	1.04408e-17
C183	A!#4	VDD#8	2.27391e-17
C184	GND#26	VDD#34	3.84815e-18
C185	VDD#39	VDD#20	1.0238e-17
C186	VDD#26	CIN#7	4.04071e-18
C187	net3#2	SOUT#6	1.96305e-17
C188	GND#32	VDD#35	1.10177e-17
C189	SOUT#10	CIN#9	4.46078e-17
C190	XI1/XI4/net24#9	XI1/XI4/net24#13	6.59037e-18
C191	net3#16	SOUT#24	5.32835e-17
C192	RST#2	GND#38	7.88615e-18
C193	A!#6	CIN#3	5.33566e-18
C194	XI1/XI4/net24#13	XI1/XI4/net24#2	1.71266e-17
C195	XI1/XI4/net24#11	SOUT#14	9.22297e-18
C196	XI1/D#19	GND#35	1.62572e-18
C197	GND#32	VDD#34	7.62525e-17
C198	PHI!#3	XI1/D	3.80638e-17
C199	SOUT#10	B!#11	3.84272e-17
C200	A!#9	CIN#3	1.29853e-18
C201	PHI#5	VDD#22	5.40385e-18
C202	COUT#6	RST#4	4.68358e-17
C203	GND#38	PHI#3	3.38517e-18
C204	VDD#8	SOUT#1	4.22292e-18
C205	PHI!#4	PHI!#5	5.34824e-18
C206	VDD#42	VDD#10	1.0238e-17
C207	SOUT#11	net3#16	1.58573e-18
C208	GND#32	VDD#27	2.62509e-18
C209	GND#4	PHI#3	5.08165e-18
C210	VDD#24	XI0/XI1/net2#3	5.00211e-18
C211	SOUT#4	CIN#4	4.68557e-18
C212	VDD#26	B!#3	8.47855e-18
C213	SOUT#14	XI1/Q	7.83548e-18
C214	VDD#22	VDD#30	7.96099e-18
C215	XI1/D#19	GND#12	2.47983e-18
C216	VDD#2	A!#4	5.50567e-17
C217	PHI!#2	XI1/XI4/net24	3.28269e-17
C218	GND#18	XI1/Q#2	5.13993e-18
C219	GND#35	XI1/D#2	5.80251e-18
C220	SOUT#11	net3#9	2.43834e-17
C221	CIN#11	RST#3	1.2685e-18
C222	B!#1	A!#3	4.63673e-17
C223	B!#10	CIN#13	8.34923e-17
C224	SOUT#6	CIN#5	3.39838e-18
C225	VDD#37	XI0/XI1/net2#3	3.05777e-18
C226	B!#14	B!#4	7.00366e-18
C227	GND#20	GND#33	8.84679e-18
C228	A!#9	CIN#2	4.96964e-17
C229	GND#12	XI1/D#2	9.24969e-18
C230	XI1/D	XI1/XI4/net24#3	2.52567e-18
C231	B!#5	SOUT#1	4.41626e-18
C232	A!#6	B!#7	5.35017e-18
C233	VDD#18	XI1/XI4/net24#11	6.3155e-17
C234	PHI#2	VDD#4	6.00445e-18
C235	SOUT#24	A!#3	2.93467e-18
C236	VDD#35	VDD	4.3302e-17
C237	A!#4	VDD#44	1.1119e-17
C238	CIN#2	A!#4	3.09365e-18
C239	RST#4	COUT#3	7.49192e-18
C240	VDD#28	VDD	5.73743e-17
C241	COUT#1	XI0/XI1/net2#3	6.65581e-18
C242	SOUT#14	SOUT#15	6.95608e-18
C243	GND#22	GND#21	7.74457e-18
C244	B!#5	CIN#13	4.0898e-17
C245	XI1/XI4/net24#13	XI1/Q#7	3.21387e-18
C246	XI1/XI4/net24#11	VDD#31	1.56401e-17
C247	GND#35	GND#34	5.35008e-18
C248	SOUT#8	A!#1	2.40961e-17
C249	XI1/XI4/net24	XI1/D#4	2.39789e-18
C250	XI0/XI1/net2#15	COUT#1	6.80992e-18
C251	B!#7	A!#9	3.9822e-18
C252	SOUT#20	XI0/XI1/net2#3	1.51276e-18
C253	A!#3	CIN#9	1.57734e-18
C254	VDD#38	XI0/XI1/net2#2	4.26212e-18
C255	VDD#27	XI1/Q	2.29012e-18
C256	PHI#5	XI1/XI4/net24	8.89281e-18
C257	VDD#42	net3#3	2.93418e-18
C258	VDD#4	VDD#33	7.96099e-18
C259	XI1/XI4/net24#3	PHI#6	4.68747e-17
C260	A!#6	SOUT#3	2.75761e-18
C261	CIN#13	VDD#16	1.37205e-17
C262	VDD#14	VDD#13	3.34678e-18
C263	VDD#10	net3#3	3.96888e-18
C264	XI1/D#17	PHI#6	1.97458e-18
C265	VDD#24	XI0/XI1/net2#2	8.46721e-18
C266	VDD#38	VDD#24	8.34952e-18
C267	GND#34	CIN#4	3.80483e-18
C268	CIN#13	VDD#42	1.34565e-17
C269	A!#9	SOUT#3	2.35212e-17
C270	XI0/XI1/net2#15	COUT#6	8.91913e-18
C271	GND#36	GND#35	9.23803e-18
C272	GND#38	GND#37	2.50799e-18
C273	SOUT#24	B!#11	2.12646e-17
C274	PHI!#6	PHI#3	9.47309e-18
C275	GND#6	CIN#3	1.73249e-18
C276	XI1/D#17	XI1/Q#12	5.0264e-17
C277	XI1/Q#12	PHI!#2	2.90831e-18
C278	XI1/Q#9	XI1/Q#11	1.53602e-18
C279	B!#10	A!#9	3.8104e-17
C280	CIN#2	SOUT#2	1.06752e-17
C281	PHI#6	XI1/Q#3	3.05252e-18
C282	XI0/XI1/net2#13	COUT#6	8.8501e-18
C283	PHI!#9	PHI#3	1.27134e-18
C284	GND#34	XI1/XI4/net24#3	4.14351e-18
C285	XI0/XI1/net2#13	GND#34	1.3169e-17
C286	XI1/Q#7	XI1/Q#5	9.68451e-18
C287	XI1/Q#6	PHI!#2	2.75539e-18
C288	GND#12	GND#16	1.79538e-17
C289	XI0/XI1/net2#16	SOUT#5	2.87586e-18
C290	GND#8	GND#37	1.02095e-17
C291	VDD#2	VDD	1.49508e-17
C292	CIN#11	VDD#42	2.19629e-17
C293	GND#16	XI1/XI4/net24#3	3.76841e-18
C294	VDD#44	VDD	4.49131e-17
C295	CIN#9	SOUT#9	3.7545e-17
C296	COUT#1	COUT#2	7.3184e-18
C297	GND#10	GND#9	7.9864e-18
C298	SOUT#14	PHI#5	1.23563e-17
C299	GND#27	SOUT#10	7.13064e-18
C300	GND#28	B!#2	3.63595e-18
C301	XI1/Q#12	XI1/D#20	2.27533e-17
C302	net3#9	VDD#39	3.67334e-17
C303	XI0/XI1/net2#13	COUT#3	3.28469e-18
C304	XI1/D#4	PHI#4	1.07136e-17
C305	GND#33	SOUT#16	1.37047e-17
C306	CIN#2	VDD#1	2.42465e-18
C307	VDD#4	VDD	1.68456e-17
C308	RST#2	net3#2	3.74826e-18
C309	VDD#33	VDD	1.01965e-16
C310	A!#9	SOUT#2	2.69483e-18
C311	A!#4	B!#10	2.23946e-18
C312	VDD#5	VDD	2.11985e-17
C313	GND#34	PHI#6	5.83194e-18
C314	RST#2	GND#34	3.10681e-18
C315	GND#22	SOUT#10	1.12163e-17
C316	GND#14	B!#2	1.48416e-18
C317	CIN#11	SOUT#6	1.79032e-18
C318	A!#4	VDD	9.31981e-18
C319	VDD#37	XI0/XI1/net2#2	1.54384e-18
C320	GND#14	GND#13	5.66199e-18
C321	GND#16	PHI#6	1.372e-18
C322	XI1/Q#11	XI1/XI4/net24#12	2.96161e-17
C323	SOUT#19	XI1/Q#2	6.59904e-18
C324	SOUT#5	RST#2	3.72778e-17
C325	GND#18	SOUT#16	4.02114e-17
C326	A!#4	SOUT#2	5.09768e-18
C327	VDD#10	CIN#11	2.53619e-17
C328	PHI!#9	VDD	4.78049e-18
C329	GND#33	SOUT#19	3.10131e-18
C330	net3#4	VDD#39	1.43985e-17
C331	PHI!#4	VDD	2.14306e-17
C332	XI1/Q#6	XI1/D#20	8.15881e-17
C333	XI1/XI4/net24#2	XI1/Q#12	1.3891e-17
C334	XI0/XI1/net2#15	SOUT#20	5.36179e-18
C335	XI1/D#10	VDD	1.26139e-17
C336	SOUT#20	RST#4	3.33183e-17
C337	PHI#5	XI1/Q	1.18127e-17
C338	VDD#41	SOUT#6	4.21273e-18
C339	VDD#8	VDD	5.6201e-18
C340	SOUT#11	B!#14	3.25292e-18
C341	VDD#43	VDD	1.8633e-17
C342	B!#11	SOUT#22	7.22189e-18
C343	VDD#26	B!#4	1.39714e-18
C344	VDD#14	VDD#18	3.92434e-17
C345	SOUT#16	SOUT#17	4.09771e-18
C346	A!#4	B!#5	1.10776e-17
C347	VDD#12	SOUT#6	4.07255e-18
C348	VDD#20	net3#4	3.89417e-17
C349	PHI!#9	PHI#2	6.19281e-17
C350	XI1/XI4/net24#6	GND#12	3.31137e-17
C351	VDD#39	XI0/XI1/net2#15	1.7071e-18
C352	B!#5	VDD	8.81226e-18
C353	XI1/XI4/net24#13	PHI#5	9.76906e-18
C354	B!#4	CIN#7	2.43471e-17
C355	XI1/Q#9	XI1/XI4/net24#3	1.58103e-18
C356	VDD#42	VDD	1.94359e-17
C357	PHI!#2	PHI#2	1.20847e-17
C358	B!#4	VDD#37	2.37247e-18
C359	VDD#10	VDD	4.30842e-18
C360	SOUT#8	VDD#16	1.33308e-17
C361	VDD#38	VDD#37	1.81893e-17
C362	B!#9	SOUT#22	1.14292e-17
C363	XI1/D#15	RST#2	4.36037e-17
C364	CIN#13	VDD	7.3798e-18
C365	GND#29	SOUT#3	5.38904e-18
C366	CIN#11	VDD	6.33291e-18
C367	PHI#5	XI1/Q#7	3.39064e-17
C368	PHI#2	PHI!#4	4.3751e-18
C369	COUT#1	XI0/XI1/net2#2	5.88268e-18
C370	GND#29	GND#6	8.36698e-18
C371	net3#2	SOUT#5	3.43763e-18
C372	SOUT#22	CIN#8	5.05993e-18
C373	VDD#43	XI1/D#10	1.29802e-17
C374	GND#14	A!#2	4.32997e-18
C375	SOUT#8	VDD#40	5.47184e-18
C376	VDD#18	VDD#17	3.34678e-18
C377	VDD#41	VDD	2.56909e-17
C378	VDD#12	VDD	4.78033e-18
C379	CIN#1	SOUT#1	3.65393e-18
C380	GND#6	SOUT#3	4.36955e-18
C381	XI1/D#2	XI1/D#17	3.60142e-18
C382	XI1/Q#9	PHI#6	4.56241e-18
C383	SOUT#18	PHI#5	1.77809e-17
C384	B!#14	SOUT#22	8.50387e-18
C385	GND#27	GND#22	9.65661e-18
C386	COUT#6	XI0/XI1/net2#2	3.27874e-18
C387	VDD#22	SOUT#14	5.47166e-17
C388	XI1/Q#7	VDD	1.11747e-17
C389	XI1/Q#11	PHI#6	1.32498e-17
C390	XI1/D#15	net3	1.96101e-17
C391	XI1/Q#5	VDD	1.57977e-17
C392	GND#8	XI1/D#14	2.67745e-17
C393	RST#3	net3#3	2.67237e-18
C394	VDD#41	VDD#40	7.78826e-18
C395	VDD#32	VDD#31	6.70431e-18
C396	B!#7	B!#8	4.0203e-18
C397	VDD#14	VDD	4.49645e-18
C398	VDD#32	VDD	8.4118e-17
C399	XI1/D#17	XI1/XI4/net24#2	6.90619e-18
C400	SOUT#14	VDD#30	1.16528e-17
C401	VDD#16	VDD	8.13251e-18
C402	XI0/XI1/net2#13	CIN#4	2.31785e-18
C403	VDD#14	XI1/XI4/net24#13	1.09794e-18
C404	VDD#40	VDD	1.44935e-17
C405	COUT#3	GND#33	1.3363e-17
C406	SOUT#18	XI1/Q#2	5.04785e-18
C407	XI1/Q#6	VDD	9.99629e-18
C408	GND#2	GND#1	2.80681e-18
C409	XI0/XI1/net2#2	SOUT#20	1.29961e-17
C410	GND#30	GND#29	2.68866e-18
C411	VDD#4	VDD#3	5.45567e-18
C412	XI0/XI1/net2#16	VDD	3.04753e-18
C413	XI1/Q#7	PHI!#1	1.21362e-17
C414	XI1/D#14	GND#37	6.93982e-18
C415	SOUT#10	SOUT#22	5.91301e-18
C416	XI1/Q#9	XI1/Q#3	2.18451e-18
C417	XI1/D#20	VDD	3.67809e-18
C418	XI1/Q#5	PHI!#1	8.79316e-18
C419	XI1/D#2	PHI!#2	1.00039e-18
C420	B!#7	SOUT#3	5.63912e-18
C421	VDD#12	VDD#11	7.9864e-18
C422	GND#38	PHI!#6	1.36671e-17
C423	RST#4	GND#20	1.13456e-17
C424	GND#34	GND#33	2.95976e-18
C425	SOUT#22	B!#4	3.05678e-18
C426	PHI!#2	XI1/XI4/net24#2	5.77081e-17
C427	VDD#31	VDD	4.74455e-17
C428	VDD#14	PHI#5	1.48609e-18
C429	VDD#39	VDD	2.30186e-17
C430	VDD#20	VDD	6.98387e-18
C431	VDD#16	VDD#15	1.68878e-17
C432	XI1/Q#7	XI1/XI4/net24	6.2497e-18
C433	PHI!#1	XI1/XI4/net24	7.48941e-17
C434	XI1/D#10	net3#2	7.8648e-18
C435	GND#30	GND#2	8.47392e-18
C436	XI1/D#19	GND#37	3.09512e-17
C437	RST#4	GND#31	1.50587e-17
C438	COUT#5	XI0/XI1/net2#2	1.85354e-18
C439	B!#10	CIN#2	2.57031e-18
C440	VDD#10	VDD#12	4.32491e-18
C441	VDD#26	VDD#37	1.09613e-17
C442	XI1/D#2	XI1/XI4/net24#2	4.04498e-17
C443	XI1/Q#5	XI1/XI4/net24	3.34152e-18
C444	XI1/XI4/net24#11	VDD	4.65294e-18
C445	VDD#24	COUT#1	5.50567e-17
C446	net3#9	VDD	1.98755e-17
C447	XI1/D#19	PHI!	3.65766e-18
C448	VDD#14	PHI!#1	3.64808e-18
C449	net3#4	VDD	2.62323e-17
C450	XI1/D#15	net3#2	3.59645e-18
C451	XI1/Q#5	VDD#14	6.35763e-17
C452	SOUT#6	CIN#6	3.8605e-18
C453	XI1/XI4/net24#4	XI1/Q#12	2.8824e-17
C454	RST#4	GND#34	3.06476e-18
C455	XI1/Q#7	VDD#32	1.95651e-18
C456	VDD#5	VDD#6	5.04192e-18
C457	VDD#32	PHI!#1	4.411e-18
C458	GND#4	PHI!#6	4.09153e-17
C459	GND#33	SOUT#18	1.33829e-17
C460	XI1/XI4/net24#6	XI1/XI4/net24#5	6.84508e-18
C461	GND#32	XI0/XI1/net2#2	1.86055e-18
C462	SOUT#7	A!#1	5.39732e-17
C463	XI0/XI1/net2#16	CIN#5	2.63779e-17
C464	CIN#11	XI1/D#14	5.73862e-18
C465	B!#11	CIN#9	3.59305e-18
C466	SOUT#24	B!#2	5.12165e-17
C467	VDD#22	VDD	6.22879e-18
C468	XI1/XI4/net24	XI1/D#3	2.28624e-18
C469	VDD#27	XI1/Q#2	2.47832e-18
C470	SOUT#5	CIN#5	4.43091e-17
C471	VDD#30	VDD	8.65204e-17
C472	GND#2	GND#6	3.86512e-18
C473	VDD#38	VDD	2.13492e-17
C474	VDD#34	XI0/XI1/net2#2	1.25381e-18
C475	GND#18	SOUT#18	3.57926e-18
C476	VDD#24	VDD	7.41165e-18
C477	VDD#14	XI1/XI4/net24	6.41722e-18
C478	A!#9	CIN#13	5.07397e-18
C479	XI1/Q#5	VDD#32	1.53345e-17
C480	VDD#32	XI1/XI4/net24	4.3074e-18
C481	VDD#26	VDD	1.04322e-17
C482	XI0/XI1/net2#16	SOUT#6	5.16806e-18
C483	VDD#37	VDD	4.07404e-17
C484	VDD#8	VDD#43	8.75267e-18
C485	VDD#22	SOUT	4.08336e-18
C486	SOUT	VDD#30	4.02348e-17
C487	SOUT#14	VDD	9.18799e-18
C488	COUT#5	RST#4	4.02246e-17
C489	XI1/D#19	PHI#3	2.62196e-18
C490	COUT#1	VDD	8.9569e-18
C491	A!#1	CIN#7	1.29274e-18
C492	XI1/D#16	XI1/D#15	9.34038e-18
C493	GND#20	COUT#3	4.01983e-17
C494	XI1/D#3	PHI#4	5.34502e-17
C495	SOUT#22	VDD	9.32721e-18
C496	VDD#20	VDD#19	8.26154e-18
C497	GND#8	GND#10	4.32491e-18
C498	GND#8	net3	4.05515e-18
C499	SOUT#20	VDD	7.57372e-18
C500	VDD#38	SOUT#20	2.939e-18
C501	SOUT#18	VDD	2.72899e-18
C502	GND#35	GND#12	1.01892e-17
C503	VDD#40	VDD#39	7.31304e-18
C504	SOUT#8	SOUT#11	8.1418e-18
C505	COUT#7	VDD	1.11412e-17
C506	COUT#5	VDD	1.10414e-17
C507	B!#2	A!#2	6.91036e-17
C508	SOUT#14	SOUT	3.34613e-17
C509	GND#26	VDD	2.72245e-17
C510	XI1/D#2	XI1/XI4/net24#4	1.54296e-18
C511	GND#37	net3	4.15538e-18
C512	GND#32	VDD	6.08273e-18
C513	SOUT#16	SOUT#19	1.38255e-17
C514	XI1/D#17	XI1/XI4/net24#4	3.52091e-17
C515	VDD#34	VDD	9.24489e-17
C516	XI1/XI4/net24#9	XI1/Q#12	4.73578e-18
C517	XI1/Q#6	PHI#5	4.16718e-17
C518	VDD#27	VDD	1.08467e-16
C519	SOUT#24	A!#2	7.14175e-18
C520	PHI#4	XI1/Q	2.93097e-18
C521	CIN#2	VDD	2.30792e-18
C522	CIN#6	XI0/XI1/net2#3	1.19235e-18
C523	GND#29	B!#7	1.31853e-17
C524	VDD#24	SOUT#20	4.20867e-18
C525	XI0/XI1/net2#13	XI0/XI1/net2	2.66668e-18
C526	PHI#2	VDD	6.79796e-17
C527	XI1/Q#6	XI1/XI4/net24	1.04447e-18
C528	XI1/XI4/net24#2	XI1/XI4/net24#4	1.52005e-18
C529	SOUT#2	VDD	9.00561e-18
C530	XI1/Q#6	VDD#31	1.9494e-18
C531	PHI#5	PHI!#2	4.78246e-17
C532	net3#2	VDD	4.21525e-17
C533	CIN#11	VDD#41	6.81056e-18
C534	XI0/XI1/net2#13	RST#2	2.21589e-17
C535	CIN#7	B!#3	5.54788e-17
C536	VDD#16	SOUT#7	8.24977e-18
C537	SOUT#11	A!#2	1.22267e-18
C538	PHI!#2	VDD	3.27746e-18
C539	GND#33	XI1/Q#3	2.16945e-18
C540	VDD#37	COUT#1	1.49363e-17
C541	RST#2	GND#8	1.03647e-17
C542	SOUT	VDD#27	1.47154e-17
C543	RST#4	XI0/XI1/net2	1.47319e-17
C544	net3#4	XI0/XI1/net2#15	3.27011e-17
C545	PHI!#6	PHI!#7	4.46757e-18
C546	B!#10	SOUT#2	7.02063e-18
C547	net3#16	B!#11	1.66613e-17
C548	GND#27	SOUT#22	9.0763e-18
C549	VDD#40	SOUT#7	2.63522e-18
C550	GND#20	SOUT#20	5.18901e-18
C551	GND#18	XI1/Q#3	4.41398e-18
C552	XI1/D#14	net3	2.44048e-18
C553	GND#34	XI1/D#17	4.75796e-18
C554	RST#2	GND#37	6.31281e-18
C555	XI1/D#4	VDD	8.75864e-18
C556	B!#5	SOUT#2	1.8238e-17
C557	PHI#5	VDD	5.43061e-17
C558	XI1/D#20	XI1/D#4	9.89326e-18
C559	GND#6	B!#7	4.04959e-17
C560	VDD#16	A!#1	4.13602e-18
C561	XI0/XI1/net2#2	VDD	5.47535e-18
C562	net3#16	B!#9	1.54183e-17
C563	CIN#11	VDD#12	1.45498e-17
C564	VDD#4	PHI!#4	5.54873e-17
C565	B!#4	VDD	1.9561e-18
C566	VDD#40	A!#1	1.82797e-18
C567	SOUT#2	VDD#42	4.81645e-18
C568	XI1/Q#12	XI1/XI4/net24#13	1.81624e-17
C569	PHI!	PHI#2	5.78599e-17
C570	VDD#26	SOUT#22	3.77905e-17
C571	GND#16	XI1/D#17	1.61841e-17
C572	GND#33	XI0/XI1/net2	2.76367e-18
C573	GND#27	CIN#9	4.17672e-18
C574	CIN#11	RST#2	7.73029e-18
C575	XI1/D#20	PHI#5	2.73964e-17
C576	net3#9	B!#9	3.8466e-18
C577	GND#22	CIN#9	2.55369e-18
C578	VDD#2	VDD#44	8.75267e-18
C579	VDD#14	XI1/D#3	1.58831e-18
C580	COUT#3	SOUT#16	2.93637e-18
C581	XI1/Q#9	GND#18	1.36992e-17
C582	COUT#3	COUT#4	4.31453e-18
C583	CIN#2	SOUT#3	2.27501e-18
C584	GND#34	XI1/XI4/net24#4	2.22377e-18
C585	XI1/D#14	RST#2	5.02859e-17
C586	PHI!#4	VDD#33	1.16528e-17
C587	B!	CIN#13	7.26056e-17
C588	VDD#42	net3#2	8.21861e-18
C589	CIN#1	VDD	2.10514e-17
C590	XI0/XI1/net2#15	SOUT#5	5.93898e-18
C591	net3#9	B!#14	1.0739e-17
C592	RST#3	VDD	2.21559e-17
C593	PHI#1	VDD	2.39701e-17
C594	A!#2	CIN#8	2.92703e-18
C595	SOUT#1	VDD	7.47753e-18
C596	GND#16	XI1/XI4/net24#4	3.29561e-18
C597	GND#32	RST#4	2.41904e-17
C598	VDD#18	XI1/XI4/net24	1.58831e-18
C599	SOUT#20	VDD#37	2.36483e-17
C600	net3#3	VDD	4.47542e-18
C601	GND#18	GND#17	2.9443e-18
C602	SOUT#6	VDD	1.22001e-17
C603	VDD#10	net3#2	1.39754e-17
C604	PHI!#1	VDD	1.47213e-17
C605	VDD#44	VDD#43	5.79597e-18
C606	GND#27	SOUT#9	2.67289e-18
C607	XI1/XI4/net24	VDD	9.38808e-18
C608	SOUT#24	B!	6.83291e-18
C609	XI0/XI1/net2#13	SOUT#5	2.17512e-17
C610	XI1/D#19	PHI!#3	2.23795e-18
C611	SOUT#7	VDD	3.25902e-18
C612	VDD#14	VDD#32	1.16687e-17
C613	GND#10	SOUT#4	4.09574e-18
C614	RST#2	net3	2.28596e-17
C615	A!#1	VDD	5.29805e-18
C616	XI1/D#14	GND#10	1.27886e-17
C617	CIN#6	VDD	1.13782e-17
C618	XI1/D#20	VDD#18	2.68757e-17
C619	GND#22	SOUT#9	5.27208e-18
C620	XI1/D#3	VDD	4.65131e-18
C621	GND#20	XI0/XI1/net2	4.49691e-18
C622	XI1/Q#7	XI1/Q#6	6.43966e-18
C623	PHI#4	VDD	5.74562e-18
C624	CIN#13	SOUT#2	6.17276e-17
C625	B!#7	A!	1.04908e-18
C626	A!	B!#10	3.24511e-17
C627	GND#28	net3#16	1.74589e-17
C628	VDD#20	XI0/XI1/net2#16	1.4293e-18
C629	CIN#7	VDD	5.19162e-18
C630	GND#36	SOUT#4	3.19662e-18
C631	CIN#13	A!	1.96333e-18
C632	XI1/D#4	PHI#5	2.70764e-17
C633	XI1/Q	VDD	2.04814e-17
C634	SOUT#16	XI1/Q#3	4.25775e-18
C635	B!#3	VDD	4.09757e-18
C636	GND#27	GND#26	2.49619e-18
C637	RST#2	SOUT#4	2.05565e-17
C638	XI0/XI1/net2#3	VDD	8.39596e-18
C639	SOUT	XI1/Q	2.45177e-18
C640	SOUT#11	A!#1	8.09714e-18
C641	XI1/D#6	XI1/D#5	4.49187e-18
C642	SOUT#19	XI1/Q#3	5.30351e-18
C643	SOUT#16	SOUT#18	1.30075e-17
C644	VDD#20	VDD#24	4.45572e-18
C645	CIN#5	XI0/XI1/net2#2	4.87283e-18
C646	XI1/D#4	VDD#18	4.83878e-18
C647	COUT#7	VDD#37	6.72863e-18
C648	XI1/D#20	VDD#31	2.76988e-18
C649	GND#22	GND#26	8.143e-18
C650	B!#2	B!	5.65793e-18
C651	VDD#41	VDD#12	1.0238e-17
C652	B!	A!#2	5.5446e-17
C653	VDD#8	B!#5	5.45177e-17
C654	B!	CIN#8	1.09996e-17
C655	SOUT#11	CIN#8	1.51494e-17
C656	RST#2	GND#10	1.18488e-17
C657	XI1/D#4	VDD#31	2.24036e-18
C658	GND#8	GND#7	7.83801e-18
C659	GND#36	PHI!#3	3.59673e-18
C660	SOUT#19	SOUT#18	3.97522e-17
C661	net3	SOUT#5	4.53739e-18
C662	XI1/Q#12	XI1/XI4/net24#12	1.90043e-17
C663	VDD#2	CIN#1	5.53658e-18
C664	XI1/XI4/net24#9	XI1/D#17	7.8821e-18
C665	VDD#34	RST#4	1.68597e-17
C666	B!#11	B!#9	1.98917e-17
C667	SOUT#22	CIN#9	1.80819e-18
C668	PHI#5	XI1/Q#2	2.86692e-17
C669	XI1/XI4/net24#9	PHI!#3	8.28164e-18
C670	VDD#39	A!#1	2.05454e-18
C671	SOUT	VDD	1.40835e-17
C672	VDD#24	VDD#23	9.27333e-18
C673	XI1/Q#9	XI1/Q#8	3.3441e-18
C674	RST#2	GND#36	9.1293e-18
C675	VDD#44	CIN#1	2.66145e-18
C676	CIN#11	net3#2	4.32779e-17
C677	XI1/XI4/net24#11	VDD#22	1.81513e-17
C678	COUT#1	SOUT#20	4.64768e-17
C679	PHI	VDD	1.81982e-17
C680	SOUT#14	SOUT#18	1.9793e-17
C681	XI1/XI4/net24#6	PHI!#3	5.17189e-18
C682	GND#36	XI1/D#19	1.4499e-17
C683	SOUT#2	VDD#41	3.04495e-18
C684	XI1/XI4/net24#6	XI1/D#17	1.49758e-18
C685	A!	B!	4.84817e-17
C686	SOUT#3	B!#2	1.91621e-18
C687	XI1/D#12	VDD#44	1.34081e-17
C688	net3#11	VDD	7.88116e-18
C689	XI0/XI1/net2#12	SOUT#5	1.10754e-18
C690	XI1/D#12	VDD	1.03077e-17
C691	GND#2	GND	2.72738e-17
C692	GND#37	GND	4.94454e-17
C693	GND#22	GND	8.80845e-18
C694	XI0/XI1/XI0/net13#2	GND#34	1.2558e-17
C695	XI0/XI1/net2#9	VDD#40	1.45156e-17
C696	GND#30	GND	5.24592e-17
C697	XI1/XI5/net13#5	RST#1	3.93763e-18
C698	GND#8	GND	6.87795e-18
C699	GND#27	GND	7.75707e-17
C700	GND#23	GND	4.72899e-17
C701	XI1/D#12	XI1/D#10	3.29649e-17
C702	net3#14	GND#27	2.13647e-17
C703	GND#31	GND	6.87042e-17
C704	XI1/XI5/net13#5	XI1/XI5/net13#3	1.64955e-17
C705	GND#20	GND	6.01736e-18
C706	net3#6	VDD	9.42787e-18
C707	GND#24	GND	4.58697e-17
C708	XI1/XI5/net13#3	XI1/XI5/net13	1.34019e-18
C709	XI0/XI1/XI0/net13#2	XI0/XI1/XI0/net13	1.47724e-18
C710	VDD#39	XI0/XI1/net2#5	7.24405e-18
C711	VDD#12	XI0/XI1/net2#9	5.4106e-17
C712	GND#14	net3#18	3.11839e-17
C713	net3#11	net3#6	4.94255e-18
C714	net3#18	B!#1	2.2742e-18
C715	XI0/XI1/net2#9	CIN#5	1.21173e-18
C716	XI1/XI5/net13#5	GND#37	2.13809e-18
C717	XI0/XI1/net2#5	VDD	4.80889e-18
C718	XI1/XI5/net13#3	RST#1	9.65375e-19
C719	XI1/D#6	XI1/XI5/net13#5	5.1354e-17
C720	VDD#16	net3#11	6.15635e-17
C721	net3#14	net3#13	4.02418e-18
C722	GND#18	GND	5.52938e-18
C723	XI1/XI5/net13#3	GND#8	5.08633e-17
C724	GND#33	GND	4.55382e-17
C725	XI0/XI1/net2#9	SOUT#6	3.59424e-18
C726	XI1/D#7	VDD#10	5.38883e-17
C727	XI0/XI1/XI0/net13#4	RST#2	1.62165e-17
C728	XI1/D#7	net3#3	3.56068e-18
C729	XI0/XI1/XI0/net13#2	GND#35	6.62433e-18
C730	CIN#8	net3#6	3.2757e-18
C731	VDD#40	XI0/XI1/net2#5	1.30927e-17
C732	XI1/D#12	XI1/D#11	2.72982e-18
C733	GND#6	GND	8.45704e-18
C734	XI0/XI1/XI0/net13#4	XI0/XI1/XI0/net13#5	1.39985e-18
C735	GND#14	GND	1.6487e-17
C736	XI1/XI5/net13#3	GND#37	1.99937e-17
C737	VDD#5	XI1/D#12	5.07001e-17
C738	XI0/XI1/net2#12	XI0/XI1/net2#13	2.34358e-17
C739	GND#29	GND	7.77858e-17
C740	GND#28	GND	1.00923e-16
C741	XI1/D#12	RST#3	3.8218e-18
C742	XI0/XI1/net2#9	VDD	5.99038e-18
C743	net3#11	A!#1	7.57752e-18
C744	VDD#43	XI1/D#7	2.1907e-17
C745	net3#18	net3#14	2.75659e-18
C746	XI1/XI5/net13#5	XI1/XI5/net13#4	1.49662e-18
C747	GND#12	GND	3.49127e-18
C748	XI1/D#12	XI1/D#7	7.31544e-18
C749	net3#11	VDD#39	1.92499e-17
C750	B!#14	net3#6	2.48359e-17
C751	net3#18	net3#16	1.59412e-17
C752	GND#35	GND	1.33841e-17
C753	XI0/XI1/net2#12	RST#2	1.33951e-17
C754	net3#18	B!#2	2.19446e-18
C755	net3#14	SOUT#10	1.90893e-17
C756	RST#2	XI1/XI5/net13#5	1.58559e-17
C757	XI0/XI1/net2#12	CIN#4	3.76602e-18
C758	GND#32	GND	6.1076e-17
C759	net3#18	SOUT#24	2.45036e-17
C760	GND#10	XI0/XI1/XI0/net13#4	5.09118e-17
C761	CIN#8	net3#11	2.44833e-18
C762	net3#6	VDD#38	2.08719e-17
C763	GND#26	GND	9.60882e-17
C764	XI1/XI5/net13#5	XI1/D#16	5.59845e-19
C765	B!#11	net3#14	4.26313e-18
C766	net3#14	GND#22	3.12965e-17
C767	XI1/D#7	XI1/D#8	2.66591e-18
C768	net3#6	B!#3	4.16658e-18
C769	net3#14	CIN#9	4.12965e-18
C770	RST#2	XI0/XI1/XI0/net13#2	1.6172e-17
C771	net3#18	GND#28	1.88957e-17
C772	XI1/D#7	VDD	1.03467e-17
C773	XI0/XI1/net2#5	net3#4	2.59209e-17
C774	XI0/XI1/net2#12	XI0/XI1/net2#10	3.45593e-18
C775	net3#6	net3#7	1.46041e-17
C776	XI0/XI1/XI0/net13#4	GND#35	1.71714e-17
C777	XI0/XI1/XI0/net13#4	XI0/XI1/XI0/net13#2	1.64955e-17
C778	net3#11	net3#10	1.44781e-17
C779	net3#14	SOUT#9	2.33071e-18
C780	XI0/XI1/net2#5	SOUT#6	1.13988e-18
C781	XI0/XI1/XI0/net13#2	XI0/XI1/net2#12	4.69308e-17
C782	XI0/XI1/net2#9	net3#4	1.93606e-17
C783	net3#18	A!#3	4.06446e-18
C784	net3#6	CIN#7	7.64271e-18
C785	XI0/XI1/net2#5	VDD#20	5.76534e-17
C786	XI0/XI1/net2#12	XI0/XI1/net2	9.43555e-19
C787	GND#36	GND	2.21981e-17
C788	SOUT#11	net3#11	2.7157e-17
C789	XI0/XI1/net2#5	CIN#6	4.5401e-18
C790	net3#6	VDD#26	6.12834e-17
C791	XI0/XI1/net2#12	GND#20	4.27062e-18
C792	GND#10	GND	5.81248e-18
C793	net3#18	net3#17	4.03534e-18
C794	GND#4	GND	2.90341e-17
C795	XI1/XI5/net13#3	RST#2	1.58114e-17
C796	net3#11	net3#9	3.21725e-17
C797	XI0/XI1/net2#9	XI0/XI1/net2#5	1.75638e-17
C798	GND#38	GND	3.20677e-17
C799	XI1/D#10	XI1/D#7	3.3989e-17
C800	net3#9	net3#6	2.46594e-17
C801	XI0/XI1/net2#12	GND#34	2.09627e-17
C802	XI1/D#15	XI1/XI5/net13#5	1.42469e-18
C803	XI1/XI5/net13#5	GND#38	1.65357e-17
C804	XI1/XI5/net13#3	XI1/D#15	1.98365e-18
C805	GND#16	GND	3.53956e-18
C806	net3#16	net3#14	1.21367e-17
C807	net3#11	SOUT#7	4.09829e-18
C808	GND#34	GND	2.93302e-17
C809	VDD#41	XI0/XI1/net2#9	6.37152e-18
C810	XI0/XI1/net2#9	XI0/XI1/net2#7	1.56189e-18
C811	XI0/XI1/net2#5	XI0/XI1/net2#4	1.50642e-18
C812	B!#14	A!#1	6.36598e-19
C813	B!#11	A!#2	7.40945e-19
C814	B!#9	A!#2	8.71941e-19
C815	CIN#13	A!#1	6.60017e-19
C816	A!#1	CIN#8	8.2626e-19
C817	B!#5	CIN#1	9.33843e-19
C818	B!#7	CIN#3	1.29331e-18
C819	GND#26	B!#3	6.89259e-19
C820	GND#26	B!#4	7.03248e-19
C821	GND#14	CIN#13	6.67183e-19
C822	GND#20	CIN#4	7.67752e-19
C823	GND#2	CIN#2	8.17588e-19
C824	GND#26	CIN#8	1.04902e-18
C825	net3#16	A!#3	5.87684e-19
C826	net3#6	A!#1	7.6486e-19
C827	SOUT#3	B!#1	7.91083e-19
C828	B!#2	SOUT#8	7.93386e-19
C829	SOUT#24	B!#1	8.11212e-19
C830	B!#5	SOUT#7	8.45903e-19
C831	B!#10	SOUT#3	9.04773e-19
C832	SOUT#22	B!#3	9.38469e-19
C833	B!#4	VDD#38	7.31422e-19
C834	VDD#37	B!#3	1.12447e-18
C835	B!#14	VDD#38	1.24021e-18
C836	CIN#1	RST#3	8.92617e-19
C837	net3#16	B!#2	6.23458e-19
C838	SOUT#24	CIN#9	5.74591e-19
C839	CIN#13	SOUT#11	8.62763e-19
C840	CIN#13	SOUT#1	9.73491e-19
C841	VDD#12	CIN#6	4.8046e-19
C842	CIN#5	VDD	5.05446e-19
C843	VDD#24	CIN#6	8.61141e-19
C844	CIN#2	VDD#8	1.30482e-18
C845	CIN#13	VDD#40	1.40846e-18
C846	net3#18	CIN#9	3.7252e-19
C847	net3#11	CIN#6	3.75673e-19
C848	net3#4	CIN#11	4.08444e-19
C849	net3#9	CIN#7	7.33206e-19
C850	net3#11	CIN#7	7.62892e-19
C851	net3#16	CIN#9	9.2752e-19
C852	XI1/D#14	CIN#4	1.47002e-18
C853	RST	GND#38	7.64175e-19
C854	GND#35	RST#2	9.48137e-19
C855	COUT#7	VDD#26	1.06668e-18
C856	GND#26	SOUT#10	5.8379e-19
C857	GND#8	SOUT#4	6.94836e-19
C858	GND#26	SOUT#9	8.94058e-19
C859	GND#14	SOUT#3	1.60329e-18
C860	SOUT#19	PHI#6	8.86585e-19
C861	XI1/D#15	GND#37	1.19132e-18
C862	XI1/D#14	GND#36	1.22071e-18
C863	COUT#5	XI0/XI1/net2	7.55169e-19
C864	GND#12	XI1/XI4/net24#3	9.20398e-19
C865	GND#12	XI1/XI4/net24#2	9.87977e-19
C866	GND#33	XI1/Q#2	4.8289e-19
C867	XI1/D#19	PHI#2	8.74572e-19
C868	XI1/XI4/net24#2	PHI#6	7.75967e-19
C869	XI1/XI4/net24#2	PHI#5	9.535e-19
C870	XI1/Q#12	PHI#5	7.94002e-19
C871	VDD#34	SOUT#20	5.92296e-19
C872	VDD#10	SOUT#6	6.94836e-19
C873	SOUT#11	VDD#39	7.64293e-19
C874	SOUT	VDD#28	7.94421e-19
C875	VDD#16	SOUT#1	1.21155e-18
C876	SOUT#11	VDD	1.24623e-18
C877	SOUT#8	VDD	2.30293e-18
C878	VDD#42	SOUT#1	2.33481e-18
C879	XI1/XI4/net24#12	PHI!#2	5.31333e-19
C880	SOUT#2	net3#3	5.53224e-19
C881	net3#2	SOUT#1	5.64483e-19
C882	net3#3	SOUT#6	9.94394e-19
C883	SOUT#1	net3#3	1.14891e-18
C884	XI1/D#14	SOUT#4	7.99321e-19
C885	XI1/D#2	SOUT#4	8.55242e-19
C886	XI1/D#15	SOUT#5	1.40543e-18
C887	VDD#41	net3#4	7.43559e-19
C888	VDD#40	net3#4	1.13006e-18
C889	SOUT#14	XI1/Q#2	9.16304e-19
C890	XI1/D#12	net3#3	5.3688e-19
C891	XI1/D#6	net3	5.92325e-19
C892	XI1/D#16	net3	6.12214e-19
C893	XI0/XI1/net2#13	SOUT#4	4.31906e-19
C894	XI0/XI1/net2#5	SOUT#7	6.36383e-19
C895	VDD#34	XI0/XI1/net2#3	6.35307e-19
C896	XI1/XI4/net24#4	XI1/D#4	6.43942e-19
C897	XI1/XI4/net24#12	XI1/D#4	7.95905e-19
C898	XI0/XI1/net2#5	net3#10	3.92263e-19
C899	XI1/D#20	XI1/Q	3.0256e-19
C900	XI1/D#17	XI1/Q#3	3.77893e-19
C901	XI1/Q#6	XI1/D#4	4.04483e-19
C902	XI1/Q#5	XI1/D#3	4.90626e-19
C903	XI1/D#17	XI1/Q#2	5.79029e-19
C904	XI1/D#4	XI1/Q	6.8315e-19
C905	XI1/XI4/net24#4	XI1/Q#2	6.00447e-19
C906	A!	GND	4.26025e-17
C907	B!	GND	1.80451e-17
C908	CIN	GND	4.37666e-17
C909	COUT	GND	5.80222e-17
C910	PHI	GND	2.63637e-17
C911	PHI!	GND	2.61452e-17
C912	RST	GND	4.74996e-17
C913	SOUT	GND	1.90083e-17
C914	VDD	GND	3.20589e-19
C915	XI0/XI0/net4	GND	3.66456e-19
C916	XI1/XI4/net9	GND	3.18655e-19
C917	XI1/XI4/net25	GND	3.17892e-19
C918	XI0/XI1/net2#3	GND	3.13736e-18
C919	B!#3	GND	1.96891e-18
C920	XI1/Q	GND	2.99886e-18
C921	CIN#7	GND	4.03466e-18
C922	PHI#4	GND	1.97867e-18
C923	XI1/D#3	GND	2.28632e-20
C924	CIN#6	GND	1.05456e-18
C925	A!#1	GND	1.42922e-17
C926	SOUT#7	GND	6.82093e-19
C927	XI1/XI4/net24	GND	4.03648e-18
C928	PHI!#1	GND	4.28642e-19
C929	SOUT#6	GND	7.98051e-18
C930	net3#3	GND	1.99398e-18
C931	SOUT#1	GND	5.3701e-19
C932	RST#3	GND	2.24078e-17
C933	CIN#1	GND	1.94181e-18
C934	XI0/XI1/net2	GND	2.79716e-17
C935	SOUT#9	GND	6.61416e-18
C936	XI1/Q#3	GND	1.48647e-17
C937	CIN#9	GND	1.2684e-17
C938	PHI#6	GND	1.79318e-17
C939	XI1/XI4/net24#3	GND	9.99763e-18
C940	CIN#4	GND	3.26818e-17
C941	A!#3	GND	1.01721e-17
C942	B!#1	GND	5.70285e-18
C943	XI1/D	GND	6.5331e-18
C944	PHI!#3	GND	1.96485e-17
C945	SOUT#4	GND	1.79942e-17
C946	net3	GND	3.35095e-17
C947	SOUT#3	GND	2.67248e-17
C948	PHI#3	GND	5.87414e-17
C949	RST#1	GND	1.1724e-17
C950	CIN#3	GND	3.0384e-17
C951	B!#4	GND	1.36471e-17
C952	SOUT#10	GND	2.85374e-17
C953	XI0/XI1/net2#2	GND	4.81417e-17
C954	XI1/Q#2	GND	5.16577e-17
C955	CIN#8	GND	5.83005e-17
C956	PHI#5	GND	5.15321e-17
C957	XI1/D#4	GND	4.17494e-19
C958	XI1/XI4/net24#4	GND	1.30667e-17
C959	CIN#5	GND	4.82674e-17
C960	A!#2	GND	4.77762e-17
C961	SOUT#8	GND	2.47467e-17
C962	B!#2	GND	2.1597e-17
C963	XI1/XI4/net24#2	GND	1.89551e-17
C964	XI1/D#2	GND	1.32495e-17
C965	PHI!#2	GND	4.45746e-17
C966	SOUT#5	GND	7.09963e-17
C967	net3#2	GND	2.87717e-17
C968	SOUT#2	GND	4.38104e-17
C969	PHI#2	GND	7.00049e-17
C970	RST#2	GND	1.11901e-16
C971	CIN#2	GND	9.12433e-17
C972	VDD#27	GND	6.12471e-17
C973	VDD#34	GND	5.19488e-17
C974	COUT#5	GND	2.86579e-17
C975	COUT#7	GND	5.5611e-17
C976	SOUT#18	GND	4.39033e-17
C977	SOUT#20	GND	6.34412e-17
C978	SOUT#22	GND	3.17079e-17
C979	COUT#3	GND	8.6743e-18
C980	COUT#6	GND	1.18843e-17
C981	COUT#1	GND	1.10825e-17
C982	SOUT#14	GND	3.23517e-18
C983	SOUT#19	GND	1.85261e-17
C984	SOUT#16	GND	8.43156e-18
C985	VDD#26	GND	3.11409e-18
C986	VDD#24	GND	2.60645e-19
C987	VDD#38	GND	2.30328e-19
C988	VDD#22	GND	2.25295e-18
C989	net3#6	GND	3.57652e-19
C990	B!#14	GND	9.80247e-18
C991	B!#9	GND	2.71264e-17
C992	B!#11	GND	1.8348e-17
C993	XI0/XI1/net2#13	GND	1.75343e-17
C994	XI0/XI1/net2#15	GND	2.92719e-17
C995	net3#4	GND	6.19466e-18
C996	net3#9	GND	7.68778e-18
C997	net3#16	GND	2.01534e-17
C998	XI1/XI4/net24#11	GND	2.17241e-18
C999	XI1/XI4/net24#12	GND	1.17061e-17
C1000	XI1/Q#11	GND	2.17936e-17
C1001	XI1/Q#9	GND	1.09498e-17
C1002	XI0/XI1/net2#12	GND	8.07284e-18
C1003	VDD#20	GND	3.74949e-19
C1004	VDD#39	GND	3.8563e-19
C1005	VDD#18	GND	1.60408e-18
C1006	SOUT#11	GND	1.47042e-17
C1007	SOUT#24	GND	1.90347e-17
C1008	XI1/D#20	GND	3.08439e-18
C1009	XI1/D#17	GND	1.03645e-17
C1010	XI0/XI1/net2#16	GND	6.12784e-18
C1011	XI1/Q#6	GND	4.30485e-18
C1012	XI1/Q#12	GND	1.07724e-17
C1013	VDD#40	GND	2.20805e-19
C1014	VDD#16	GND	1.74351e-18
C1015	VDD#32	GND	2.81797e-20
C1016	VDD#14	GND	6.91838e-19
C1017	XI0/XI1/XI0/net13#4	GND	1.30885e-17
C1018	XI0/XI1/net2#9	GND	6.73319e-19
C1019	XI1/Q#5	GND	2.09121e-18
C1020	XI1/Q#7	GND	2.16707e-19
C1021	XI1/XI4/net24#13	GND	1.93822e-17
C1022	XI1/XI4/net24#6	GND	7.33202e-18
C1023	XI1/XI4/net24#9	GND	1.65682e-17
C1024	VDD#12	GND	6.90231e-19
C1025	XI1/D#19	GND	3.40898e-17
C1026	XI1/D#14	GND	2.50795e-17
C1027	CIN#11	GND	2.54598e-17
C1028	CIN#13	GND	4.20471e-17
C1029	VDD#10	GND	4.14886e-19
C1030	B!#5	GND	1.84278e-19
C1031	B!#10	GND	1.80502e-17
C1032	B!#7	GND	2.11962e-17
C1033	XI1/D#7	GND	8.64157e-19
C1034	XI1/XI5/net13#3	GND	1.06358e-17
C1035	VDD#43	GND	1.23303e-18
C1036	VDD#8	GND	2.68286e-19
C1037	XI1/D#15	GND	3.82381e-17
C1038	XI1/D#10	GND	6.97924e-18
C1039	PHI!#4	GND	1.77609e-18
C1040	PHI!#9	GND	3.36789e-17
C1041	PHI!#6	GND	2.42088e-17
C1042	A!#4	GND	9.82776e-18
C1043	A!#9	GND	3.5289e-17
C1044	A!#6	GND	1.02907e-17
C1045	VDD#5	GND	3.60805e-19
C1046	VDD#4	GND	1.26825e-18
C1047	XI1/D#6	GND	1.74398e-17
C1048	XI1/D#16	GND	2.47453e-17
C1049	VDD#44	GND	7.14874e-20
C1050	VDD#2	GND	8.37146e-19
C1051	VDD#25	GND	3.24858e-19
C1052	VDD#7	GND	1.61383e-19
C1053	XI1/Q#8	GND	8.40992e-20
C1054	XI1/XI5/net13#5	GND	1.07127e-17
C1055	XI1/D#12	GND	5.19077e-18
C1056	XI0/XI1/XI0/net13#2	GND	1.40813e-17
C1057	XI0/XI1/net2#5	GND	1.61789e-18
C1058	net3#11	GND	3.5721e-19
C1059	net3#14	GND	8.13405e-18
C1060	net3#18	GND	6.35766e-18
C1061	PHI#7	GND	5.02545e-17
C1062	RST#4	GND	9.43711e-17
*
*
.ENDS HA_ACCUM
*
