** Post-Layout Supply Voltage Characterization
** Sweeping Vdd from 0.85V to 1.10V

** Include model files
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45n1svt.inc'
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45p1svt.inc'
.include 'NAND_X1-post-layout.sp'

** Parameter definition for sweep
.param supply=1.0

.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0
+    POST=1

** Power supplies
Vgnd gnd 0 0
Vsupply vdd 0 supply

** Input stimulus that scales with supply voltage
** Input A: transitions for measuring tpdr and tpdf
Va a 0 PWL(0n 0 0.5n 0 0.51n supply 1.0n supply 1.01n 0 1.5n 0 1.51n supply 2.0n supply)

** Input B: held high
Vb b 0 supply

** Instantiate the extracted cell
** Port order from .SUBCKT: A B GND VDD Y
Xnand a b gnd vdd y NAND_X1

** Load capacitance
Cload y 0 5e-15

** Transient analysis with parameter sweep
.tran 1p 2n SWEEP supply 0.85 1.10 0.05

** Measurements for tpdr (falling A, rising Y)
.MEASURE TRAN tpdr
+ TRIG=v(a) VAL='0.5*supply' FALL=1
+ TARG=v(y) VAL='0.5*supply' RISE=1

** Measurements for tpdf (rising A, falling Y)
.MEASURE TRAN tpdf
+ TRIG=v(a) VAL='0.5*supply' RISE=1
+ TARG=v(y) VAL='0.5*supply' FALL=1

** Rise time measurement for input A
.MEASURE TRAN tr_a
+ TRIG=v(a) VAL='0.1*supply' RISE=1
+ TARG=v(a) VAL='0.9*supply' RISE=1

** Fall time measurement for input A  
.MEASURE TRAN tf_a
+ TRIG=v(a) VAL='0.9*supply' FALL=1
+ TARG=v(a) VAL='0.1*supply' FALL=1

** Rise time measurement for output Y
.MEASURE TRAN tr_y
+ TRIG=v(y) VAL='0.2*supply' RISE=1
+ TARG=v(y) VAL='0.8*supply' RISE=1

** Fall time measurement for output Y
.MEASURE TRAN tf_y
+ TRIG=v(y) VAL='0.8*supply' FALL=1
+ TARG=v(y) VAL='0.2*supply' FALL=1

** Static current measurement (when output is stable high, beginning of simulation)
.MEASURE TRAN istat AVG I(Vsupply) FROM=50p TO=150p

** Peak current measurement
.MEASURE TRAN ipeak MIN I(Vsupply) FROM=0p TO=2n

** Print statements for waveform viewing
.print tran v(a) v(b) v(y) i(Vsupply)

.END
