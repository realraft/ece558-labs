** Half Adder Accumulator SPICE Netlist with Testbench
** step3_zguro_raftery.sp

** Parameter for clock period
.param tclk=1n

** Temperature and Options
.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0
+    POST=1
+    PROBE=1

** Include GPDK045 transistor models
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45n1svt.inc'
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45p1svt.inc'

** Library name: components
** Cell name: INV
** View name: schematic
.subckt INV a gnd vdd y
mpm0 y a vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm0 y a gnd gnd g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9
.ends INV

** Library name: components
** Cell name: XOR
** View name: schematic
.subckt XOR a b gnd vdd y
mpm3 y a net11 vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mpm2 net11 net9 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mpm1 y net5 net4 vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mpm0 net4 b vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mnm3 net18 b gnd gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm2 net15 net9 gnd gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm1 y a net18 gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm0 y net5 net15 gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
xi1 b gnd vdd net9 INV
xi0 a gnd vdd net5 INV
.ends XOR

** Library name: components
** Cell name: NAND
** View name: schematic
.subckt NAND a b gnd vdd y
mpm1 y a vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mpm0 y b vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm1 net13 b gnd gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm0 y a net13 gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
.ends NAND

** Library name: components
** Cell name: AND
** View name: schematic
.subckt AND a b gnd vdd y
xi0 a b gnd vdd net2 NAND
xi2 net2 gnd vdd y INV
.ends AND

** Library name: components
** Cell name: HA
** View name: schematic
.subckt HA a b c gnd s vdd
xi0 a b gnd vdd s XOR
xi1 a b gnd vdd c AND
.ends HA

** Library name: components
** Cell name: RST-FF
** View name: schematic
.subckt RST_FF gnd phi rst s sout vdd
mpm3 net14 net6 net11 vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mpm2 net11 net7 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mpm1 net7 phi net4 vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mpm0 net4 net5 vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6
mnm3 net22 net7 net19 gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm2 net14 phi net22 gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm1 net15 net5 net19 gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
mnm0 net7 net6 net15 gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9
xi1 phi gnd vdd net6 INV
xi0 net14 gnd vdd sout INV
xi2 rst s gnd vdd net5 NAND
.ends RST_FF

** Main Circuit: HA_ACCUM
** Top level subcircuit
.subckt HA_ACCUM cin phi rst cout sout gnd vdd
xi0 cin sout cout gnd net3 vdd HA
xi1 gnd phi rst net3 sout vdd RST_FF
.ends HA_ACCUM

** Test Circuit Instantiation
xdut cin phi rst cout sout 0 vdd HA_ACCUM

** Power Supply - NO vgnd LINE!
vvdd vdd 0 DC 1.1

** Load capacitances on outputs
Ccout cout 0 5f
Csout sout 0 5f

** Include vector file for stimulus
.vec 'step3_zguro_raftery.vec'

** Transient Analysis
.tran 1p 6n

** Measurements for propagation delays and rise/fall times
** Measure propagation delays (50% to 50%)
.measure tran tpdr_sout trig v(phi) val=0.55 rise=2 
+                       targ v(sout) val=0.55 rise=1
.measure tran tpdf_sout trig v(phi) val=0.55 rise=3 
+                       targ v(sout) val=0.55 fall=1

.measure tran tpdr_cout trig v(phi) val=0.55 rise=4 
+                       targ v(cout) val=0.55 rise=1
.measure tran tpdf_cout trig v(phi) val=0.55 rise=4 
+                       targ v(cout) val=0.55 fall=1

** Measure rise and fall times (20% to 80%)
.measure tran tr_sout trig v(sout) val=0.22 rise=1 
+                     targ v(sout) val=0.88 rise=1
.measure tran tf_sout trig v(sout) val=0.88 fall=1 
+                     targ v(sout) val=0.22 fall=1

.measure tran tr_cout trig v(cout) val=0.22 rise=1 
+                     targ v(cout) val=0.88 rise=1
.measure tran tf_cout trig v(cout) val=0.88 fall=1 
+                     targ v(cout) val=0.22 fall=1

** Print statements for debugging
.print tran v(phi) v(rst) v(cin) v(sout) v(cout)

.END
