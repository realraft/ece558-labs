** Generated for: hspiceD
** Generated on: Sep 30 20:03:28 2025
** Design library name: NAND_X1
** Design cell name: NAND_X1
** Design view name: schematic

** Model includes
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45n1svt.inc'
.include '/opt/cadence/gpdk045/gpdk045_v_6_0/models/hspice/g45p1svt.inc'


.param vdd_val=1.1

.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0

.vec 'input.vec'

** Power supplies with current measurement
Vgnd gnd 0 0

Vsupply vdd 0 vdd_val

** Library name: NAND_X1
** Cell name: NAND_X1
** View name: schematic
mpm1 y a vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm0 y b vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm1 net13 b gnd gnd g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm0 y a net13 net13 g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1

Cload y 0 5e-15

** Transient analysis
.tran 1p 2.5n

** HSPICE Delay Measurements
** Propagation delay rising (tpdr) - when A falls, Y rises
.MEASURE TRAN tpdr
+ TRIG=v(a) VAL='0.5*vdd_val' FALL=1
+ TARG=v(y) VAL='0.5*vdd_val' RISE=1

** Propagation delay falling (tpdf) - when A rises, Y falls
.MEASURE TRAN tpdf
+ TRIG=v(a) VAL='0.5*vdd_val' RISE=1
+ TARG=v(y) VAL='0.5*vdd_val' FALL=1

** Rise time of output Y (tr) - 20%-80% metric
.MEASURE TRAN tr_y
+ TRIG=v(y) VAL='0.2*vdd_val' RISE=1
+ TARG=v(y) VAL='0.8*vdd_val' RISE=1

** Fall time of output Y (tf) - 80%-20% metric
.MEASURE TRAN tf_y
+ TRIG=v(y) VAL='0.8*vdd_val' FALL=1
+ TARG=v(y) VAL='0.2*vdd_val' FALL=1

** Static leakage current measurement (when both inputs are low - first vector)
.MEASURE TRAN istat AVG I(Vsupply) FROM=50p TO=150p

** Peak current measurement during entire simulation
.MEASURE TRAN ipeak MIN I(Vsupply) FROM=0p TO=2.5n

.print tran v(a) v(b) v(y) i(Vsupply)
.option post

.END
