*
*
*
*                       LINUX           Tue Nov 11 21:24:14 2025
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 24.1.0-p089
*  Build Date     : Wed Dec 18 09:06:09 PST 2024
*
*  HSPICE LIBRARY
*
*  QRC_TECH_DIR /ece558_658/pdk/verification/qrc/typical 
*
*
*

*
.SUBCKT 4BIT_ACCUM CIN COUT GND PHI RST SOUT0 SOUT1 SOUT2 SOUT3 VDD
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MXI3/XI0/XI0/XI1/MNM0	XI3/XI0/XI0/BNOT#8	SOUT3#3	GND#71	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI3/XI1/XI5/MNM1	XI3/XI1/XI5/net13	XI3/net1	GND#73	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI0/XI1/XI0/MNM1	XI3/XI0/XI1/XI0/net13#5	SOUT3#4	GND#75
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI1/XI4/MNM0	XI3/XI1/XI4/net24#5	XI3/XI1/XI4/PHINOT#3
+ XI3/XI1/XI4/net36	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI1/XI4/MNM3	XI3/XI1/XI4/net36	XI3/XI1/D	GND#77	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI0/XI0/MNM2	XI3/XI0/XI0/net15	XI3/XI0/XI0/BNOT	GND#79
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI3/XI0/XI0/MNM0	XI3/net1#17	XI3/XI0/XI0/ANOT#3
+ XI3/XI0/XI0/net15	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI3/XI0/XI1/XI0/MNM0	XI3/XI0/XI1/net2#10	net21#4
+ XI3/XI0/XI1/XI0/net13	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI1/XI4/MNM2	XI3/XI1/XI4/net25	XI3/XI1/XI4/net24#3	GND#81
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI1/XI4/MNM1	XI3/XI1/Q#8	PHI#24	XI3/XI1/XI4/net25	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI0/XI0/MNM1	XI3/net1#13	net21#9	XI3/XI0/XI0/net18
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI3/XI1/XI6/MNM0	SOUT3#17	XI3/XI1/Q#3	GND#83	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI3/XI0/XI0/MNM3	XI3/XI0/XI0/net18	SOUT3#9	GND#87	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI3/XI0/XI1/XI2/MNM0	COUT#4	XI3/XI0/XI1/net2	GND#85	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI2/XI0/XI0/XI1/MNM0	XI2/XI0/XI0/BNOT#8	SOUT2#3	GND#49	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI2/XI1/XI5/MNM1	XI2/XI1/XI5/net13	XI2/net1	GND#51	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI0/XI1/XI0/MNM1	XI2/XI0/XI1/XI0/net13#5	SOUT2#4	GND#53
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI1/XI4/MNM0	XI2/XI1/XI4/net24#5	XI2/XI1/XI4/PHINOT#3
+ XI2/XI1/XI4/net36	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI1/XI4/MNM3	XI2/XI1/XI4/net36	XI2/XI1/D	GND#55	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI0/XI0/MNM2	XI2/XI0/XI0/net15	XI2/XI0/XI0/BNOT	GND#57
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI2/XI0/XI0/MNM0	XI2/net1#17	XI2/XI0/XI0/ANOT#3
+ XI2/XI0/XI0/net15	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI2/XI0/XI1/XI0/MNM0	XI2/XI0/XI1/net2#10	net14#4
+ XI2/XI0/XI1/XI0/net13	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI1/XI4/MNM2	XI2/XI1/XI4/net25	XI2/XI1/XI4/net24#3	GND#59
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI1/XI4/MNM1	XI2/XI1/Q#8	PHI#18	XI2/XI1/XI4/net25	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI0/XI0/MNM1	XI2/net1#13	net14#9	XI2/XI0/XI0/net18
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI2/XI1/XI6/MNM0	SOUT2#17	XI2/XI1/Q#3	GND#61	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI2/XI0/XI0/MNM3	XI2/XI0/XI0/net18	SOUT2#9	GND#65	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI2/XI0/XI1/XI2/MNM0	net21#13	XI2/XI0/XI1/net2	GND#63	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI1/XI0/XI0/XI1/MNM0	XI1/XI0/XI0/BNOT#8	SOUT1#3	GND#27	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI1/XI1/XI5/MNM1	XI1/XI1/XI5/net13	XI1/net1	GND#29	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI0/XI1/XI0/MNM1	XI1/XI0/XI1/XI0/net13#5	SOUT1#4	GND#31
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI1/XI4/MNM0	XI1/XI1/XI4/net24#5	XI1/XI1/XI4/PHINOT#3
+ XI1/XI1/XI4/net36	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI1/XI4/MNM3	XI1/XI1/XI4/net36	XI1/XI1/D	GND#33	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI0/XI0/MNM2	XI1/XI0/XI0/net15	XI1/XI0/XI0/BNOT	GND#35
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI1/XI0/XI0/MNM0	XI1/net1#17	XI1/XI0/XI0/ANOT#3
+ XI1/XI0/XI0/net15	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI1/XI0/XI1/XI0/MNM0	XI1/XI0/XI1/net2#10	net7#4	XI1/XI0/XI1/XI0/net13
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI1/XI4/MNM2	XI1/XI1/XI4/net25	XI1/XI1/XI4/net24#3	GND#37
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI1/XI4/MNM1	XI1/XI1/Q#8	PHI#12	XI1/XI1/XI4/net25	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI0/XI0/MNM1	XI1/net1#13	net7#9	XI1/XI0/XI0/net18	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI1/XI1/XI6/MNM0	SOUT1#17	XI1/XI1/Q#3	GND#39	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI1/XI0/XI0/MNM3	XI1/XI0/XI0/net18	SOUT1#9	GND#43	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI1/XI0/XI1/XI2/MNM0	net14#13	XI1/XI0/XI1/net2	GND#41	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI0/XI0/XI0/XI1/MNM0	XI0/XI0/XI0/BNOT#8	SOUT0#3	GND#5	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI0/XI1/XI5/MNM1	XI0/XI1/XI5/net13	XI0/net1	GND#7	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI0/XI1/XI0/MNM1	XI0/XI0/XI1/XI0/net13#5	SOUT0#4	GND#9
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI1/XI4/MNM0	XI0/XI1/XI4/net24#5	XI0/XI1/XI4/PHINOT#3
+ XI0/XI1/XI4/net36	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI1/XI4/MNM3	XI0/XI1/XI4/net36	XI0/XI1/D	GND#11	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI0/XI0/MNM2	XI0/XI0/XI0/net15	XI0/XI0/XI0/BNOT	GND#13
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI0/XI0/XI0/MNM0	XI0/net1#17	XI0/XI0/XI0/ANOT#3
+ XI0/XI0/XI0/net15	GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI0/XI0/XI1/XI0/MNM0	XI0/XI0/XI1/net2#10	CIN#4	XI0/XI0/XI1/XI0/net13
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI1/XI4/MNM2	XI0/XI1/XI4/net25	XI0/XI1/XI4/net24#3	GND#15
+ GND	g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI1/XI4/MNM1	XI0/XI1/Q#8	PHI#6	XI0/XI1/XI4/net25	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI0/XI0/XI0/MNM1	XI0/net1#13	CIN#9	XI0/XI0/XI0/net18	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=1.44e-14	PD=7.6e-07	PS=6e-07
+ sa=1.4e-07 sb=2.45e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI0/XI1/XI6/MNM0	SOUT0#17	XI0/XI1/Q#3	GND#17	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI0/XI0/XI0/MNM3	XI0/XI0/XI0/net18	SOUT0#9	GND#21	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=1.44e-14	AS=3.36e-14	PD=6e-07	PS=7.6e-07
+ sa=2.45e-07 sb=1.4e-07 sca=5.51597 scb=0.00169014 scc=6.16736e-06 fw=2.4e-07
MXI0/XI0/XI1/XI2/MNM0	net7#13	XI0/XI0/XI1/net2	GND#19	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI0/XI0/XI0/XI0/MNM0	XI0/XI0/XI0/ANOT#7	CIN#3	GND#1	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.90867 scb=0.00164474 scc=3.75172e-06 fw=1.2e-07
MXI0/XI1/XI5/MNM0	XI0/XI1/D#5	RST#1	XI0/XI1/XI5/net13#4	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.82604 scb=0.000193838 scc=1.85478e-08 fw=2.4e-07
MXI0/XI1/XI4/XI1/MNM0	XI0/XI1/XI4/PHINOT#7	PHI#3	GND#3	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.99885 scb=0.00021225 scc=1.92763e-08 fw=1.2e-07
MXI1/XI0/XI0/XI0/MNM0	XI1/XI0/XI0/ANOT#7	net7#3	GND#23	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI1/XI1/XI5/MNM0	XI1/XI1/D#5	RST#4	XI1/XI1/XI5/net13#4	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI1/XI1/XI4/XI1/MNM0	XI1/XI1/XI4/PHINOT#7	PHI#9	GND#25	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI2/XI0/XI0/XI0/MNM0	XI2/XI0/XI0/ANOT#7	net14#3	GND#45	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI2/XI1/XI5/MNM0	XI2/XI1/D#5	RST#7	XI2/XI1/XI5/net13#4	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI2/XI1/XI4/XI1/MNM0	XI2/XI1/XI4/PHINOT#7	PHI#15	GND#47	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI3/XI0/XI0/XI0/MNM0	XI3/XI0/XI0/ANOT#7	net21#3	GND#67	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.52044 scb=0.00152619 scc=3.72446e-06 fw=1.2e-07
MXI3/XI1/XI5/MNM0	XI3/XI1/D#5	RST#10	XI3/XI1/XI5/net13#4	GND
+ g45n1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MXI3/XI1/XI4/XI1/MNM0	XI3/XI1/XI4/PHINOT#7	PHI#21	GND#69	GND
+ g45n1svt	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MXI3/XI0/XI0/XI1/MPM0	XI3/XI0/XI0/BNOT#6	SOUT3#1	VDD#85	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI3/XI1/XI5/MPM0	XI3/XI1/D#8	XI3/net1#3	VDD#87	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI3/XI0/XI1/XI0/MPM0	XI3/XI0/XI1/net2#7	SOUT3#6	VDD#89	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI3/XI1/XI4/MPM3	XI3/XI1/Q#4	XI3/XI1/XI4/PHINOT
+ XI3/XI1/XI4/net17	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI3/XI1/XI4/MPM2	XI3/XI1/XI4/net17	XI3/XI1/XI4/net24	VDD#91
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI3/XI0/XI0/MPM0	XI3/XI0/XI0/net4	SOUT3#7	VDD#93	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI3/XI0/XI0/MPM1	XI3/net1#10	XI3/XI0/XI0/ANOT
+ XI3/XI0/XI0/net4	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI3/XI0/XI1/XI0/MPM1	XI3/XI0/XI1/net2#4	net21#6	VDD#97	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI3/XI1/XI4/MPM0	XI3/XI1/XI4/net9	XI3/XI1/D#3	VDD#95	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI3/XI1/XI4/MPM1	XI3/XI1/XI4/net24#10	PHI#22	XI3/XI1/XI4/net9
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI3/XI0/XI0/MPM3	XI3/net1#7	net21#7	XI3/XI0/XI0/net11
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI3/XI1/XI6/MPM0	SOUT3#15	XI3/XI1/Q	VDD#99	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
MXI3/XI0/XI0/MPM2	XI3/XI0/XI0/net11	XI3/XI0/XI0/BNOT#3	VDD#103
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI3/XI0/XI1/XI2/MPM0	COUT#2	XI3/XI0/XI1/net2#3	VDD#101	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 fw=2.4e-07
MXI2/XI0/XI0/XI1/MPM0	XI2/XI0/XI0/BNOT#6	SOUT2#1	VDD#59	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI2/XI1/XI5/MPM0	XI2/XI1/D#8	XI2/net1#3	VDD#61	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI2/XI0/XI1/XI0/MPM0	XI2/XI0/XI1/net2#7	SOUT2#6	VDD#63	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI2/XI1/XI4/MPM3	XI2/XI1/Q#4	XI2/XI1/XI4/PHINOT
+ XI2/XI1/XI4/net17	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI2/XI1/XI4/MPM2	XI2/XI1/XI4/net17	XI2/XI1/XI4/net24	VDD#65
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI2/XI0/XI0/MPM0	XI2/XI0/XI0/net4	SOUT2#7	VDD#67	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI2/XI0/XI0/MPM1	XI2/net1#10	XI2/XI0/XI0/ANOT
+ XI2/XI0/XI0/net4	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI2/XI0/XI1/XI0/MPM1	XI2/XI0/XI1/net2#4	net14#6	VDD#71	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI2/XI1/XI4/MPM0	XI2/XI1/XI4/net9	XI2/XI1/D#3	VDD#69	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI2/XI1/XI4/MPM1	XI2/XI1/XI4/net24#10	PHI#16	XI2/XI1/XI4/net9
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI2/XI0/XI0/MPM3	XI2/net1#7	net14#7	XI2/XI0/XI0/net11
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI2/XI1/XI6/MPM0	SOUT2#15	XI2/XI1/Q	VDD#73	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
MXI2/XI0/XI0/MPM2	XI2/XI0/XI0/net11	XI2/XI0/XI0/BNOT#3	VDD#77
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI2/XI0/XI1/XI2/MPM0	net21#11	XI2/XI0/XI1/net2#3	VDD#75	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 fw=2.4e-07
MXI1/XI0/XI0/XI1/MPM0	XI1/XI0/XI0/BNOT#6	SOUT1#1	VDD#33	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI1/XI1/XI5/MPM0	XI1/XI1/D#8	XI1/net1#3	VDD#35	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI1/XI0/XI1/XI0/MPM0	XI1/XI0/XI1/net2#7	SOUT1#6	VDD#37	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI1/XI1/XI4/MPM3	XI1/XI1/Q#4	XI1/XI1/XI4/PHINOT
+ XI1/XI1/XI4/net17	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI1/XI1/XI4/MPM2	XI1/XI1/XI4/net17	XI1/XI1/XI4/net24	VDD#39
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI1/XI0/XI0/MPM0	XI1/XI0/XI0/net4	SOUT1#7	VDD#41	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI1/XI0/XI0/MPM1	XI1/net1#10	XI1/XI0/XI0/ANOT
+ XI1/XI0/XI0/net4	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI1/XI0/XI1/XI0/MPM1	XI1/XI0/XI1/net2#4	net7#6	VDD#45	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI1/XI1/XI4/MPM0	XI1/XI1/XI4/net9	XI1/XI1/D#3	VDD#43	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI1/XI1/XI4/MPM1	XI1/XI1/XI4/net24#10	PHI#10	XI1/XI1/XI4/net9
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI1/XI0/XI0/MPM3	XI1/net1#7	net7#7	XI1/XI0/XI0/net11	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI1/XI1/XI6/MPM0	SOUT1#15	XI1/XI1/Q	VDD#47	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
MXI1/XI0/XI0/MPM2	XI1/XI0/XI0/net11	XI1/XI0/XI0/BNOT#3	VDD#51
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI1/XI0/XI1/XI2/MPM0	net14#11	XI1/XI0/XI1/net2#3	VDD#49	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 fw=2.4e-07
MXI0/XI0/XI0/XI1/MPM0	XI0/XI0/XI0/BNOT#6	SOUT0#1	VDD#7	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI0/XI1/XI5/MPM0	XI0/XI1/D#8	XI0/net1#3	VDD#9	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI0/XI0/XI1/XI0/MPM0	XI0/XI0/XI1/net2#7	SOUT0#6	VDD#11	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI0/XI1/XI4/MPM3	XI0/XI1/Q#4	XI0/XI1/XI4/PHINOT
+ XI0/XI1/XI4/net17	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI0/XI1/XI4/MPM2	XI0/XI1/XI4/net17	XI0/XI1/XI4/net24	VDD#13
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI0/XI0/XI0/MPM0	XI0/XI0/XI0/net4	SOUT0#7	VDD#15	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI0/XI0/XI0/MPM1	XI0/net1#10	XI0/XI0/XI0/ANOT
+ XI0/XI0/XI0/net4	VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI0/XI0/XI1/XI0/MPM1	XI0/XI0/XI1/net2#4	CIN#6	VDD#19	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI0/XI1/XI4/MPM0	XI0/XI1/XI4/net9	XI0/XI1/D#3	VDD#17	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=1.4e-07 sb=2.45e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI0/XI1/XI4/MPM1	XI0/XI1/XI4/net24#10	PHI#4	XI0/XI1/XI4/net9
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=2.45e-07 sb=1.4e-07 sca=7.67082 scb=0.00406069 scc=4.89818e-05 fw=4.8e-07
MXI0/XI0/XI0/MPM3	XI0/net1#7	CIN#7	XI0/XI0/XI0/net11	VDD
+ g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=2.88e-14	PD=1.24e-06	PS=1.08e-06
+ sa=1.4e-07 sb=2.45e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI0/XI1/XI6/MPM0	SOUT0#15	XI0/XI1/Q	VDD#21	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
MXI0/XI0/XI0/MPM2	XI0/XI0/XI0/net11	XI0/XI0/XI0/BNOT#3	VDD#25
+ VDD	g45p1svt	L=4.5e-08	W=4.8e-07
+ AD=2.88e-14	AS=6.72e-14	PD=1.08e-06	PS=1.24e-06
+ sa=2.45e-07 sb=1.4e-07 sca=15.1999 scb=0.012812 scc=0.00139229 fw=4.8e-07
MXI0/XI0/XI1/XI2/MPM0	net7#11	XI0/XI0/XI1/net2#3	VDD#23	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 fw=2.4e-07
MXI0/XI0/XI0/XI0/MPM0	XI0/XI0/XI0/ANOT#5	CIN#1	VDD#1	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.95118 scb=0.00508612 scc=7.502e-05 fw=2.4e-07
MXI0/XI1/XI5/MPM1	XI0/XI1/D#11	RST#3	VDD#6	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.26407 scb=0.00404065 scc=4.42753e-05 fw=2.4e-07
MXI0/XI1/XI4/XI1/MPM0	XI0/XI1/XI4/PHINOT#5	PHI#1	VDD#3	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.1139 scb=0.00244911 scc=5.96896e-06 fw=2.4e-07
MXI1/XI0/XI0/XI0/MPM0	XI1/XI0/XI0/ANOT#5	net7	VDD#27	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI1/XI1/XI5/MPM1	XI1/XI1/D#11	RST#6	VDD#32	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI1/XI1/XI4/XI1/MPM0	XI1/XI1/XI4/PHINOT#5	PHI#7	VDD#29	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
MXI2/XI0/XI0/XI0/MPM0	XI2/XI0/XI0/ANOT#5	net14	VDD#53	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI2/XI1/XI5/MPM1	XI2/XI1/D#11	RST#9	VDD#58	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI2/XI1/XI4/XI1/MPM0	XI2/XI1/XI4/PHINOT#5	PHI#13	VDD#55	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
MXI3/XI0/XI0/XI0/MPM0	XI3/XI0/XI0/ANOT#5	net21	VDD#79	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 fw=2.4e-07
MXI3/XI1/XI5/MPM1	XI3/XI1/D#11	RST#12	VDD#84	VDD	g45p1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96481 scb=0.00395847 scc=4.42604e-05 fw=2.4e-07
MXI3/XI1/XI4/XI1/MPM0	XI3/XI1/XI4/PHINOT#5	PHI#19	VDD#81	VDD
+ g45p1svt	L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.81464 scb=0.00236693 scc=5.95408e-06 fw=2.4e-07
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rl1	CIN#1	CIN#2	306.867249	$poly_conn
Rl2	CIN#2	CIN#3	383.790314	$poly_conn
Rl3	RST#1	RST#2	76.098015	$poly_conn
Rl4	RST#2	RST#3	606.867249	$poly_conn
Rl5	PHI#1	PHI#2	199.979935	$poly_conn
Rl6	PHI#2	PHI#3	492.287628	$poly_conn
Rl7	SOUT0#1	SOUT0#2	142.287613	$poly_conn
Rl8	SOUT0#2	SOUT0#3	549.979919	$poly_conn
Rl9	XI0/net1	XI0/net1#2	622.251892	$poly_conn
Rl10	XI0/net1#2	XI0/net1#3	60.713398	$poly_conn
Rl11	SOUT0#4	SOUT0#5	215.364548	$poly_conn
Rl12	SOUT0#5	SOUT0#6	469.210693	$poly_conn
Rl13	XI0/XI1/XI4/PHINOT	XI0/XI1/XI4/PHINOT#2	206.461472
+ $poly_conn
Rl14	XI0/XI1/XI4/PHINOT#2	XI0/XI1/XI4/PHINOT#3	391.076874
+ $poly_conn
Rl15	XI0/XI1/XI4/net24	XI0/XI1/XI4/net24#2	490.321899
+ $poly_conn
Rl16	XI0/XI1/D	XI0/XI1/D#2	117.244949	$poly_conn
Rl17	SOUT0#7	SOUT0#8	101.860336	$poly_conn
Rl18	XI0/XI0/XI0/BNOT	XI0/XI0/XI0/BNOT#2	141.475723
+ $poly_conn
Rl19	XI0/XI0/XI0/ANOT	XI0/XI0/XI0/ANOT#2	372.251862
+ $poly_conn
Rl20	XI0/XI0/XI0/ANOT#2	XI0/XI0/XI0/ANOT#3	210.713394
+ $poly_conn
Rl21	CIN#4	CIN#5	418.405701	$poly_conn
Rl22	CIN#5	CIN#6	264.559540	$poly_conn
Rl23	XI0/XI1/D#3	XI0/XI1/D#4	53.014187	$poly_conn
Rl24	XI0/XI1/XI4/net24#3	XI0/XI1/XI4/net24#4	145.321869
+ $poly_conn
Rl25	PHI#4	PHI#5	126.098015	$poly_conn
Rl26	PHI#5	PHI#6	464.559570	$poly_conn
Rl27	CIN#7	CIN#8	222.251862	$poly_conn
Rl28	CIN#8	CIN#9	360.713379	$poly_conn
Rl29	XI0/XI1/Q	XI0/XI1/Q#2	449.174927	$poly_conn
Rl30	XI0/XI1/Q#2	XI0/XI1/Q#3	241.482620	$poly_conn
Rl31	XI0/XI0/XI1/net2	XI0/XI0/XI1/net2#2	560.713379
+ $poly_conn
Rl32	XI0/XI0/XI1/net2#2	XI0/XI0/XI1/net2#3	129.944168
+ $poly_conn
Rl33	XI0/XI0/XI0/BNOT#3	XI0/XI0/XI0/BNOT#4	60.706493
+ $poly_conn
Rl34	SOUT0#9	SOUT0#10	113.398796	$poly_conn
Rl35	net7	net7#2	306.867249	$poly_conn
Rl36	net7#2	net7#3	383.790314	$poly_conn
Rl37	RST#4	RST#5	76.098015	$poly_conn
Rl38	RST#5	RST#6	606.867249	$poly_conn
Rl39	PHI#7	PHI#8	199.979935	$poly_conn
Rl40	PHI#8	PHI#9	492.287628	$poly_conn
Rl41	SOUT1#1	SOUT1#2	142.287613	$poly_conn
Rl42	SOUT1#2	SOUT1#3	549.979919	$poly_conn
Rl43	XI1/net1	XI1/net1#2	622.251892	$poly_conn
Rl44	XI1/net1#2	XI1/net1#3	60.713398	$poly_conn
Rl45	SOUT1#4	SOUT1#5	215.364548	$poly_conn
Rl46	SOUT1#5	SOUT1#6	469.210693	$poly_conn
Rl47	XI1/XI1/XI4/PHINOT	XI1/XI1/XI4/PHINOT#2	206.461472
+ $poly_conn
Rl48	XI1/XI1/XI4/PHINOT#2	XI1/XI1/XI4/PHINOT#3	391.076874
+ $poly_conn
Rl49	XI1/XI1/XI4/net24	XI1/XI1/XI4/net24#2	490.321899
+ $poly_conn
Rl50	XI1/XI1/D	XI1/XI1/D#2	117.244949	$poly_conn
Rl51	SOUT1#7	SOUT1#8	101.860336	$poly_conn
Rl52	XI1/XI0/XI0/BNOT	XI1/XI0/XI0/BNOT#2	141.475723
+ $poly_conn
Rl53	XI1/XI0/XI0/ANOT	XI1/XI0/XI0/ANOT#2	372.251862
+ $poly_conn
Rl54	XI1/XI0/XI0/ANOT#2	XI1/XI0/XI0/ANOT#3	210.713394
+ $poly_conn
Rl55	net7#4	net7#5	418.405701	$poly_conn
Rl56	net7#5	net7#6	264.559540	$poly_conn
Rl57	XI1/XI1/D#3	XI1/XI1/D#4	53.014187	$poly_conn
Rl58	XI1/XI1/XI4/net24#3	XI1/XI1/XI4/net24#4	145.321869
+ $poly_conn
Rl59	PHI#10	PHI#11	126.098015	$poly_conn
Rl60	PHI#11	PHI#12	464.559570	$poly_conn
Rl61	net7#7	net7#8	222.251862	$poly_conn
Rl62	net7#8	net7#9	360.713379	$poly_conn
Rl63	XI1/XI1/Q	XI1/XI1/Q#2	449.174927	$poly_conn
Rl64	XI1/XI1/Q#2	XI1/XI1/Q#3	241.482620	$poly_conn
Rl65	XI1/XI0/XI1/net2	XI1/XI0/XI1/net2#2	560.713379
+ $poly_conn
Rl66	XI1/XI0/XI1/net2#2	XI1/XI0/XI1/net2#3	129.944168
+ $poly_conn
Rl67	XI1/XI0/XI0/BNOT#3	XI1/XI0/XI0/BNOT#4	60.706493
+ $poly_conn
Rl68	SOUT1#9	SOUT1#10	113.398796	$poly_conn
Rl69	net14	net14#2	306.867249	$poly_conn
Rl70	net14#2	net14#3	383.790314	$poly_conn
Rl71	RST#7	RST#8	76.098015	$poly_conn
Rl72	RST#8	RST#9	606.867249	$poly_conn
Rl73	PHI#13	PHI#14	199.979935	$poly_conn
Rl74	PHI#14	PHI#15	492.287628	$poly_conn
Rl75	SOUT2#1	SOUT2#2	142.287613	$poly_conn
Rl76	SOUT2#2	SOUT2#3	549.979919	$poly_conn
Rl77	XI2/net1	XI2/net1#2	622.251892	$poly_conn
Rl78	XI2/net1#2	XI2/net1#3	60.713398	$poly_conn
Rl79	SOUT2#4	SOUT2#5	215.364548	$poly_conn
Rl80	SOUT2#5	SOUT2#6	469.210693	$poly_conn
Rl81	XI2/XI1/XI4/PHINOT	XI2/XI1/XI4/PHINOT#2	206.461472
+ $poly_conn
Rl82	XI2/XI1/XI4/PHINOT#2	XI2/XI1/XI4/PHINOT#3	391.076874
+ $poly_conn
Rl83	XI2/XI1/XI4/net24	XI2/XI1/XI4/net24#2	490.321899
+ $poly_conn
Rl84	XI2/XI1/D	XI2/XI1/D#2	117.244949	$poly_conn
Rl85	SOUT2#7	SOUT2#8	101.860336	$poly_conn
Rl86	XI2/XI0/XI0/BNOT	XI2/XI0/XI0/BNOT#2	141.475723
+ $poly_conn
Rl87	XI2/XI0/XI0/ANOT	XI2/XI0/XI0/ANOT#2	372.251862
+ $poly_conn
Rl88	XI2/XI0/XI0/ANOT#2	XI2/XI0/XI0/ANOT#3	210.713394
+ $poly_conn
Rl89	net14#4	net14#5	418.405701	$poly_conn
Rl90	net14#5	net14#6	264.559540	$poly_conn
Rl91	XI2/XI1/D#3	XI2/XI1/D#4	53.014187	$poly_conn
Rl92	XI2/XI1/XI4/net24#3	XI2/XI1/XI4/net24#4	145.321869
+ $poly_conn
Rl93	PHI#16	PHI#17	126.098015	$poly_conn
Rl94	PHI#17	PHI#18	464.559570	$poly_conn
Rl95	net14#7	net14#8	222.251862	$poly_conn
Rl96	net14#8	net14#9	360.713379	$poly_conn
Rl97	XI2/XI1/Q	XI2/XI1/Q#2	449.174927	$poly_conn
Rl98	XI2/XI1/Q#2	XI2/XI1/Q#3	241.482620	$poly_conn
Rl99	XI2/XI0/XI1/net2	XI2/XI0/XI1/net2#2	560.713379
+ $poly_conn
Rl100	XI2/XI0/XI1/net2#2	XI2/XI0/XI1/net2#3	129.944168
+ $poly_conn
Rl101	XI2/XI0/XI0/BNOT#3	XI2/XI0/XI0/BNOT#4	60.706493
+ $poly_conn
Rl102	SOUT2#9	SOUT2#10	113.398796	$poly_conn
Rl103	net21	net21#2	306.867249	$poly_conn
Rl104	net21#2	net21#3	383.790314	$poly_conn
Rl105	RST#10	RST#11	76.098015	$poly_conn
Rl106	RST#11	RST#12	606.867249	$poly_conn
Rl107	PHI#19	PHI#20	199.979935	$poly_conn
Rl108	PHI#20	PHI#21	492.287628	$poly_conn
Rl109	SOUT3#1	SOUT3#2	142.287613	$poly_conn
Rl110	SOUT3#2	SOUT3#3	549.979919	$poly_conn
Rl111	XI3/net1	XI3/net1#2	622.251892	$poly_conn
Rl112	XI3/net1#2	XI3/net1#3	60.713398	$poly_conn
Rl113	SOUT3#4	SOUT3#5	215.364548	$poly_conn
Rl114	SOUT3#5	SOUT3#6	469.210693	$poly_conn
Rl115	XI3/XI1/XI4/PHINOT	XI3/XI1/XI4/PHINOT#2	206.461472
+ $poly_conn
Rl116	XI3/XI1/XI4/PHINOT#2	XI3/XI1/XI4/PHINOT#3	391.076874
+ $poly_conn
Rl117	XI3/XI1/XI4/net24	XI3/XI1/XI4/net24#2	490.321899
+ $poly_conn
Rl118	XI3/XI1/D	XI3/XI1/D#2	117.244949	$poly_conn
Rl119	SOUT3#7	SOUT3#8	101.860336	$poly_conn
Rl120	XI3/XI0/XI0/BNOT	XI3/XI0/XI0/BNOT#2	141.475723
+ $poly_conn
Rl121	XI3/XI0/XI0/ANOT	XI3/XI0/XI0/ANOT#2	372.251862
+ $poly_conn
Rl122	XI3/XI0/XI0/ANOT#2	XI3/XI0/XI0/ANOT#3	210.713394
+ $poly_conn
Rl123	net21#4	net21#5	418.405701	$poly_conn
Rl124	net21#5	net21#6	264.559540	$poly_conn
Rl125	XI3/XI1/D#3	XI3/XI1/D#4	53.014187	$poly_conn
Rl126	XI3/XI1/XI4/net24#3	XI3/XI1/XI4/net24#4	145.321869
+ $poly_conn
Rl127	PHI#22	PHI#23	126.098015	$poly_conn
Rl128	PHI#23	PHI#24	464.559570	$poly_conn
Rl129	net21#7	net21#8	222.251862	$poly_conn
Rl130	net21#8	net21#9	360.713379	$poly_conn
Rl131	XI3/XI1/Q	XI3/XI1/Q#2	449.174927	$poly_conn
Rl132	XI3/XI1/Q#2	XI3/XI1/Q#3	241.482620	$poly_conn
Rl133	XI3/XI0/XI1/net2	XI3/XI0/XI1/net2#2	560.713379
+ $poly_conn
Rl134	XI3/XI0/XI1/net2#2	XI3/XI0/XI1/net2#3	129.944168
+ $poly_conn
Rl135	XI3/XI0/XI0/BNOT#3	XI3/XI0/XI0/BNOT#4	60.706493
+ $poly_conn
Rl136	SOUT3#9	SOUT3#10	113.398796	$poly_conn
Rk1	VDD#1	VDD#2	31.000000	$metal1_conn
Rk2	GND#1	GND#2	75.000000	$metal1_conn
Rk3	XI0/XI1/D#5	XI0/XI1/D#6	37.501156	$metal1_conn
Rk4	VDD#3	VDD#4	31.000000	$metal1_conn
Rk5	VDD#5	VDD#6	31.001158	$metal1_conn
Rk6	GND#3	GND#4	75.000000	$metal1_conn
Rk7	XI0/XI0/XI0/ANOT#4	XI0/XI0/XI0/ANOT#5	31.001158
+ $metal1_conn
Rk8	XI0/XI0/XI0/ANOT#6	XI0/XI0/XI0/ANOT#7	75.001549
+ $metal1_conn
Rk9	XI0/XI1/XI4/PHINOT#4	XI0/XI1/XI4/PHINOT#5	31.001158
+ $metal1_conn
Rk10	XI0/XI1/XI4/PHINOT#6	XI0/XI1/XI4/PHINOT#7	75.001549
+ $metal1_conn
Rk11	VDD#7	VDD#8	31.000000	$metal1_conn
Rk12	XI0/XI1/XI5/net13#2	XI0/XI1/XI5/net13#3	0.001157
+ $metal1_conn
Rk13	XI0/XI1/XI5/net13#3	XI0/XI1/XI5/net13#5	0.232308
+ $metal1_conn
Rk15	XI0/XI1/XI5/net13	XI0/XI1/XI5/net13#2	37.500000
+ $metal1_conn
Rk16	XI0/XI1/XI5/net13#4	XI0/XI1/XI5/net13#5	37.500000
+ $metal1_conn
Rk17	GND#5	GND#6	75.000000	$metal1_conn
Rk18	XI0/XI1/D#7	XI0/XI1/D#9	0.001157	$metal1_conn
Rk19	XI0/XI1/D#9	XI0/XI1/D#10	0.120231	$metal1_conn
Rk20	XI0/XI1/D#10	XI0/XI1/D#12	0.114924	$metal1_conn
Rk22	XI0/XI1/D#8	XI0/XI1/D#9	31.000000	$metal1_conn
Rk23	XI0/XI1/D#11	XI0/XI1/D#12	31.000000	$metal1_conn
Rk24	XI0/XI0/XI0/BNOT#5	XI0/XI0/XI0/BNOT#6	31.001158
+ $metal1_conn
Rk25	GND#7	GND#8	37.500000	$metal1_conn
Rk26	VDD#9	VDD#10	31.000000	$metal1_conn
Rk27	XI0/XI0/XI0/BNOT#7	XI0/XI0/XI0/BNOT#8	75.001549
+ $metal1_conn
Rk28	XI0/XI1/D#14	XI0/XI1/D#15	0.450092	$metal1_conn
Rk29	XI0/XI1/D#15	XI0/XI1/D#16	0.266916	$metal1_conn
Rk30	GND#9	GND#10	37.500000	$metal1_conn
Rk31	VDD#11	VDD#12	31.000000	$metal1_conn
Rk32	XI0/XI1/Q#4	XI0/XI1/Q#5	15.500000	$metal1_conn
Rk33	XI0/XI1/XI4/net24#5	XI0/XI1/XI4/net24#6	37.500000
+ $metal1_conn
Rk34	XI0/XI1/XI4/PHINOT#2	XI0/XI1/XI4/PHINOT#9	46.516312
+ $metal1_conn
Rk35	VDD#13	VDD#14	15.500000	$metal1_conn
Rk36	GND#11	GND#12	37.500000	$metal1_conn
Rk37	VDD#15	VDD#16	15.500000	$metal1_conn
Rk38	GND#13	GND#14	37.500000	$metal1_conn
Rk39	XI0/XI1/Q#6	XI0/XI1/Q#7	0.365328	$metal1_conn
Rk40	XI0/XI0/XI0/ANOT#2	XI0/XI0/XI0/ANOT#9	46.855549
+ $metal1_conn
Rk42	XI0/XI0/XI1/XI0/net13#2	XI0/XI0/XI1/XI0/net13#4
+ 0.232308	$metal1_conn
Rk43	XI0/XI0/XI1/XI0/net13#4	XI0/XI0/XI1/XI0/net13#5
+ 37.501156	$metal1_conn
Rk44	XI0/XI0/XI1/XI0/net13	XI0/XI0/XI1/XI0/net13#2	37.500000
+ $metal1_conn
Rk46	XI0/XI0/XI1/net2#5	XI0/XI0/XI1/net2#8	0.237615
+ $metal1_conn
Rk47	XI0/XI0/XI1/net2#8	XI0/XI0/XI1/net2#9	0.001157
+ $metal1_conn
Rk48	XI0/XI0/XI1/net2#4	XI0/XI0/XI1/net2#5	31.000000
+ $metal1_conn
Rk49	XI0/XI0/XI1/net2#7	XI0/XI0/XI1/net2#8	31.000000
+ $metal1_conn
Rk50	XI0/XI1/D#17	XI0/XI1/D#2	0.292025	$metal1_conn
Rk51	XI0/XI1/D#2	XI0/XI1/D#19	0.466581	$metal1_conn
Rk52	CIN#5	CIN#11	45.731133	$metal1_conn
Rk53	SOUT0#11	SOUT0#8	0.156463	$metal1_conn
Rk54	SOUT0#8	SOUT0#2	45.836899	$metal1_conn
Rk55	VDD#17	VDD#18	15.500000	$metal1_conn
Rk56	GND#15	GND#16	37.500000	$metal1_conn
Rk57	VDD#19	VDD#20	31.001158	$metal1_conn
Rk58	XI0/XI1/XI4/net24#4	XI0/XI1/XI4/net24#2	45.402275
+ $metal1_conn
Rk59	XI0/XI1/XI4/net24#2	XI0/XI1/XI4/net24#9	0.668824
+ $metal1_conn
Rk60	XI0/XI1/D#20	XI0/XI1/D#4	45.082287	$metal1_conn
Rk61	XI0/XI1/XI4/net24#10	XI0/XI1/XI4/net24#11	15.500000
+ $metal1_conn
Rk62	XI0/XI1/XI4/net24#12	XI0/XI1/XI4/net24#13	0.688239
+ $metal1_conn
Rk63	XI0/XI1/Q#8	XI0/XI1/Q#9	37.500000	$metal1_conn
Rk64	XI0/XI0/XI1/net2#11	XI0/XI0/XI1/net2#12	0.001157
+ $metal1_conn
Rk65	XI0/XI0/XI1/net2#12	XI0/XI0/XI1/net2#13	0.169876
+ $metal1_conn
Rk66	XI0/XI0/XI1/net2#10	XI0/XI0/XI1/net2#11	37.500000
+ $metal1_conn
Rk67	XI0/net1#4	XI0/net1#2	46.295746	$metal1_conn
Rk68	XI0/XI0/XI0/BNOT#9	XI0/XI0/XI0/BNOT#10	2.761596
+ $metal1_conn
Rk69	XI0/XI0/XI0/BNOT#11	XI0/XI0/XI0/BNOT#2	45.782852
+ $metal1_conn
Rk71	XI0/net1#6	XI0/net1#9	0.322022	$metal1_conn
Rk72	XI0/net1#9	XI0/net1#11	0.257371	$metal1_conn
Rk74	XI0/net1#7	XI0/net1#6	15.500000	$metal1_conn
Rk75	XI0/net1#10	XI0/net1#11	15.500000	$metal1_conn
Rk77	XI0/net1#14	XI0/net1#16	0.305642	$metal1_conn
Rk78	XI0/net1#16	XI0/net1#18	0.240992	$metal1_conn
Rk80	XI0/net1#13	XI0/net1#14	37.500000	$metal1_conn
Rk81	XI0/net1#17	XI0/net1#18	37.500000	$metal1_conn
Rk82	CIN	CIN#12	0.221625	$metal1_conn
Rk83	CIN#12	CIN#13	0.688033	$metal1_conn
Rk84	CIN#13	CIN#8	46.508373	$metal1_conn
Rk85	VDD#21	VDD#22	31.000000	$metal1_conn
Rk86	VDD#23	VDD#24	31.000000	$metal1_conn
Rk87	GND#17	GND#18	75.000000	$metal1_conn
Rk88	GND#19	GND#20	75.000000	$metal1_conn
Rk89	XI0/XI1/Q#2	XI0/XI1/Q#11	45.453136	$metal1_conn
Rk90	XI0/XI1/Q#11	XI0/XI1/Q#12	0.376483	$metal1_conn
Rk91	XI0/XI0/XI1/net2#2	XI0/XI0/XI1/net2#15	45.440205
+ $metal1_conn
Rk92	XI0/XI0/XI1/net2#15	XI0/XI0/XI1/net2#16	0.343778
+ $metal1_conn
Rk93	XI0/XI0/XI0/BNOT#4	XI0/XI0/XI0/BNOT#14	45.156464
+ $metal1_conn
Rk94	SOUT0#14	SOUT0#15	31.001158	$metal1_conn
Rk95	VDD#25	VDD#26	15.500000	$metal1_conn
Rk96	GND#21	GND#22	37.500000	$metal1_conn
Rk97	net7#10	net7#11	31.001158	$metal1_conn
Rk98	SOUT0#16	SOUT0#17	75.001549	$metal1_conn
Rk99	net7#12	net7#13	75.001549	$metal1_conn
Rk100	SOUT0#18	SOUT0#19	1.205139	$metal1_conn
Rk101	SOUT0#20	SOUT0#5	46.880508	$metal1_conn
Rk102	SOUT0#22	SOUT0#10	0.248977	$metal1_conn
Rk103	SOUT0#10	SOUT0#24	0.776813	$metal1_conn
Rk104	net7#14	net7#15	0.885980	$metal1_conn
Rk105	VDD#27	VDD#28	31.000000	$metal1_conn
Rk106	GND#23	GND#24	75.000000	$metal1_conn
Rk107	XI1/XI1/D#5	XI1/XI1/D#6	37.501156	$metal1_conn
Rk108	VDD#29	VDD#30	31.000000	$metal1_conn
Rk109	VDD#31	VDD#32	31.001158	$metal1_conn
Rk110	GND#25	GND#26	75.000000	$metal1_conn
Rk111	XI1/XI0/XI0/ANOT#4	XI1/XI0/XI0/ANOT#5	31.001158
+ $metal1_conn
Rk112	XI1/XI0/XI0/ANOT#6	XI1/XI0/XI0/ANOT#7	75.001549
+ $metal1_conn
Rk113	XI1/XI1/XI4/PHINOT#4	XI1/XI1/XI4/PHINOT#5	31.001158
+ $metal1_conn
Rk114	XI1/XI1/XI4/PHINOT#6	XI1/XI1/XI4/PHINOT#7	75.001549
+ $metal1_conn
Rk115	VDD#33	VDD#34	31.000000	$metal1_conn
Rk116	XI1/XI1/XI5/net13#2	XI1/XI1/XI5/net13#3	0.001157
+ $metal1_conn
Rk117	XI1/XI1/XI5/net13#3	XI1/XI1/XI5/net13#5	0.232308
+ $metal1_conn
Rk119	XI1/XI1/XI5/net13	XI1/XI1/XI5/net13#2	37.500000
+ $metal1_conn
Rk120	XI1/XI1/XI5/net13#4	XI1/XI1/XI5/net13#5	37.500000
+ $metal1_conn
Rk121	GND#27	GND#28	75.000000	$metal1_conn
Rk122	XI1/XI1/D#7	XI1/XI1/D#9	0.001157	$metal1_conn
Rk123	XI1/XI1/D#9	XI1/XI1/D#10	0.120231	$metal1_conn
Rk124	XI1/XI1/D#10	XI1/XI1/D#12	0.114924	$metal1_conn
Rk126	XI1/XI1/D#8	XI1/XI1/D#9	31.000000	$metal1_conn
Rk127	XI1/XI1/D#11	XI1/XI1/D#12	31.000000	$metal1_conn
Rk128	XI1/XI0/XI0/BNOT#5	XI1/XI0/XI0/BNOT#6	31.001158
+ $metal1_conn
Rk129	GND#29	GND#30	37.500000	$metal1_conn
Rk130	VDD#35	VDD#36	31.000000	$metal1_conn
Rk131	XI1/XI0/XI0/BNOT#7	XI1/XI0/XI0/BNOT#8	75.001549
+ $metal1_conn
Rk132	XI1/XI1/D#14	XI1/XI1/D#15	0.450092	$metal1_conn
Rk133	XI1/XI1/D#15	XI1/XI1/D#16	0.266916	$metal1_conn
Rk134	GND#31	GND#32	37.500000	$metal1_conn
Rk135	VDD#37	VDD#38	31.000000	$metal1_conn
Rk136	XI1/XI1/Q#4	XI1/XI1/Q#5	15.500000	$metal1_conn
Rk137	XI1/XI1/XI4/net24#5	XI1/XI1/XI4/net24#6	37.500000
+ $metal1_conn
Rk138	XI1/XI1/XI4/PHINOT#2	XI1/XI1/XI4/PHINOT#9	46.516312
+ $metal1_conn
Rk139	VDD#39	VDD#40	15.500000	$metal1_conn
Rk140	GND#33	GND#34	37.500000	$metal1_conn
Rk141	VDD#41	VDD#42	15.500000	$metal1_conn
Rk142	GND#35	GND#36	37.500000	$metal1_conn
Rk143	XI1/XI1/Q#6	XI1/XI1/Q#7	0.365328	$metal1_conn
Rk144	XI1/XI0/XI0/ANOT#2	XI1/XI0/XI0/ANOT#9	46.855549
+ $metal1_conn
Rk146	XI1/XI0/XI1/XI0/net13#2	XI1/XI0/XI1/XI0/net13#4
+ 0.232308	$metal1_conn
Rk147	XI1/XI0/XI1/XI0/net13#4	XI1/XI0/XI1/XI0/net13#5
+ 37.501156	$metal1_conn
Rk148	XI1/XI0/XI1/XI0/net13	XI1/XI0/XI1/XI0/net13#2	37.500000
+ $metal1_conn
Rk150	XI1/XI0/XI1/net2#5	XI1/XI0/XI1/net2#8	0.237615
+ $metal1_conn
Rk151	XI1/XI0/XI1/net2#8	XI1/XI0/XI1/net2#9	0.001157
+ $metal1_conn
Rk152	XI1/XI0/XI1/net2#4	XI1/XI0/XI1/net2#5	31.000000
+ $metal1_conn
Rk153	XI1/XI0/XI1/net2#7	XI1/XI0/XI1/net2#8	31.000000
+ $metal1_conn
Rk154	XI1/XI1/D#17	XI1/XI1/D#2	0.292025	$metal1_conn
Rk155	XI1/XI1/D#2	XI1/XI1/D#19	0.466581	$metal1_conn
Rk156	net7#5	net7#17	45.731133	$metal1_conn
Rk157	SOUT1#11	SOUT1#8	0.156463	$metal1_conn
Rk158	SOUT1#8	SOUT1#2	45.836899	$metal1_conn
Rk159	VDD#43	VDD#44	15.500000	$metal1_conn
Rk160	GND#37	GND#38	37.500000	$metal1_conn
Rk161	VDD#45	VDD#46	31.001158	$metal1_conn
Rk162	XI1/XI1/XI4/net24#4	XI1/XI1/XI4/net24#2	45.402275
+ $metal1_conn
Rk163	XI1/XI1/XI4/net24#2	XI1/XI1/XI4/net24#9	0.668824
+ $metal1_conn
Rk164	XI1/XI1/D#20	XI1/XI1/D#4	45.082287	$metal1_conn
Rk165	XI1/XI1/XI4/net24#10	XI1/XI1/XI4/net24#11	15.500000
+ $metal1_conn
Rk166	XI1/XI1/XI4/net24#12	XI1/XI1/XI4/net24#13	0.688239
+ $metal1_conn
Rk167	XI1/XI1/Q#8	XI1/XI1/Q#9	37.500000	$metal1_conn
Rk168	XI1/XI0/XI1/net2#11	XI1/XI0/XI1/net2#12	0.001157
+ $metal1_conn
Rk169	XI1/XI0/XI1/net2#12	XI1/XI0/XI1/net2#13	0.169876
+ $metal1_conn
Rk170	XI1/XI0/XI1/net2#10	XI1/XI0/XI1/net2#11	37.500000
+ $metal1_conn
Rk171	XI1/net1#4	XI1/net1#2	46.295746	$metal1_conn
Rk172	XI1/XI0/XI0/BNOT#9	XI1/XI0/XI0/BNOT#10	2.761596
+ $metal1_conn
Rk173	XI1/XI0/XI0/BNOT#11	XI1/XI0/XI0/BNOT#2	45.782852
+ $metal1_conn
Rk175	XI1/net1#6	XI1/net1#9	0.322022	$metal1_conn
Rk176	XI1/net1#9	XI1/net1#11	0.257371	$metal1_conn
Rk178	XI1/net1#7	XI1/net1#6	15.500000	$metal1_conn
Rk179	XI1/net1#10	XI1/net1#11	15.500000	$metal1_conn
Rk181	XI1/net1#14	XI1/net1#16	0.305642	$metal1_conn
Rk182	XI1/net1#16	XI1/net1#18	0.240992	$metal1_conn
Rk184	XI1/net1#13	XI1/net1#14	37.500000	$metal1_conn
Rk185	XI1/net1#17	XI1/net1#18	37.500000	$metal1_conn
Rk186	net7#8	net7#19	46.508373	$metal1_conn
Rk187	net7#19	net7#20	0.688033	$metal1_conn
Rk188	net7#20	net7#21	1.364706	$metal1_conn
Rk189	VDD#47	VDD#48	31.000000	$metal1_conn
Rk190	VDD#49	VDD#50	31.000000	$metal1_conn
Rk191	GND#39	GND#40	75.000000	$metal1_conn
Rk192	GND#41	GND#42	75.000000	$metal1_conn
Rk193	XI1/XI1/Q#2	XI1/XI1/Q#11	45.453136	$metal1_conn
Rk194	XI1/XI1/Q#11	XI1/XI1/Q#12	0.376483	$metal1_conn
Rk195	XI1/XI0/XI1/net2#2	XI1/XI0/XI1/net2#15	45.440205
+ $metal1_conn
Rk196	XI1/XI0/XI1/net2#15	XI1/XI0/XI1/net2#16	0.343778
+ $metal1_conn
Rk197	XI1/XI0/XI0/BNOT#4	XI1/XI0/XI0/BNOT#14	45.156464
+ $metal1_conn
Rk198	SOUT1#14	SOUT1#15	31.001158	$metal1_conn
Rk199	VDD#51	VDD#52	15.500000	$metal1_conn
Rk200	GND#43	GND#44	37.500000	$metal1_conn
Rk201	net14#10	net14#11	31.001158	$metal1_conn
Rk202	SOUT1#16	SOUT1#17	75.001549	$metal1_conn
Rk203	net14#12	net14#13	75.001549	$metal1_conn
Rk204	SOUT1#18	SOUT1#19	1.205139	$metal1_conn
Rk205	SOUT1#20	SOUT1#5	46.880508	$metal1_conn
Rk206	SOUT1#22	SOUT1#10	0.248977	$metal1_conn
Rk207	SOUT1#10	SOUT1#24	0.776813	$metal1_conn
Rk208	net14#14	net14#15	0.885980	$metal1_conn
Rk209	VDD#53	VDD#54	31.000000	$metal1_conn
Rk210	GND#45	GND#46	75.000000	$metal1_conn
Rk211	XI2/XI1/D#5	XI2/XI1/D#6	37.501156	$metal1_conn
Rk212	VDD#55	VDD#56	31.000000	$metal1_conn
Rk213	VDD#57	VDD#58	31.001158	$metal1_conn
Rk214	GND#47	GND#48	75.000000	$metal1_conn
Rk215	XI2/XI0/XI0/ANOT#4	XI2/XI0/XI0/ANOT#5	31.001158
+ $metal1_conn
Rk216	XI2/XI0/XI0/ANOT#6	XI2/XI0/XI0/ANOT#7	75.001549
+ $metal1_conn
Rk217	XI2/XI1/XI4/PHINOT#4	XI2/XI1/XI4/PHINOT#5	31.001158
+ $metal1_conn
Rk218	XI2/XI1/XI4/PHINOT#6	XI2/XI1/XI4/PHINOT#7	75.001549
+ $metal1_conn
Rk219	VDD#59	VDD#60	31.000000	$metal1_conn
Rk220	XI2/XI1/XI5/net13#2	XI2/XI1/XI5/net13#3	0.001157
+ $metal1_conn
Rk221	XI2/XI1/XI5/net13#3	XI2/XI1/XI5/net13#5	0.232308
+ $metal1_conn
Rk223	XI2/XI1/XI5/net13	XI2/XI1/XI5/net13#2	37.500000
+ $metal1_conn
Rk224	XI2/XI1/XI5/net13#4	XI2/XI1/XI5/net13#5	37.500000
+ $metal1_conn
Rk225	GND#49	GND#50	75.000000	$metal1_conn
Rk226	XI2/XI1/D#7	XI2/XI1/D#9	0.001157	$metal1_conn
Rk227	XI2/XI1/D#9	XI2/XI1/D#10	0.120231	$metal1_conn
Rk228	XI2/XI1/D#10	XI2/XI1/D#12	0.114924	$metal1_conn
Rk230	XI2/XI1/D#8	XI2/XI1/D#9	31.000000	$metal1_conn
Rk231	XI2/XI1/D#11	XI2/XI1/D#12	31.000000	$metal1_conn
Rk232	XI2/XI0/XI0/BNOT#5	XI2/XI0/XI0/BNOT#6	31.001158
+ $metal1_conn
Rk233	GND#51	GND#52	37.500000	$metal1_conn
Rk234	VDD#61	VDD#62	31.000000	$metal1_conn
Rk235	XI2/XI0/XI0/BNOT#7	XI2/XI0/XI0/BNOT#8	75.001549
+ $metal1_conn
Rk236	XI2/XI1/D#14	XI2/XI1/D#15	0.450092	$metal1_conn
Rk237	XI2/XI1/D#15	XI2/XI1/D#16	0.266916	$metal1_conn
Rk238	GND#53	GND#54	37.500000	$metal1_conn
Rk239	VDD#63	VDD#64	31.000000	$metal1_conn
Rk240	XI2/XI1/Q#4	XI2/XI1/Q#5	15.500000	$metal1_conn
Rk241	XI2/XI1/XI4/net24#5	XI2/XI1/XI4/net24#6	37.500000
+ $metal1_conn
Rk242	XI2/XI1/XI4/PHINOT#2	XI2/XI1/XI4/PHINOT#9	46.516312
+ $metal1_conn
Rk243	VDD#65	VDD#66	15.500000	$metal1_conn
Rk244	GND#55	GND#56	37.500000	$metal1_conn
Rk245	VDD#67	VDD#68	15.500000	$metal1_conn
Rk246	GND#57	GND#58	37.500000	$metal1_conn
Rk247	XI2/XI1/Q#6	XI2/XI1/Q#7	0.365328	$metal1_conn
Rk248	XI2/XI0/XI0/ANOT#2	XI2/XI0/XI0/ANOT#9	46.855549
+ $metal1_conn
Rk250	XI2/XI0/XI1/XI0/net13#2	XI2/XI0/XI1/XI0/net13#4
+ 0.232308	$metal1_conn
Rk251	XI2/XI0/XI1/XI0/net13#4	XI2/XI0/XI1/XI0/net13#5
+ 37.501156	$metal1_conn
Rk252	XI2/XI0/XI1/XI0/net13	XI2/XI0/XI1/XI0/net13#2	37.500000
+ $metal1_conn
Rk254	XI2/XI0/XI1/net2#5	XI2/XI0/XI1/net2#8	0.237615
+ $metal1_conn
Rk255	XI2/XI0/XI1/net2#8	XI2/XI0/XI1/net2#9	0.001157
+ $metal1_conn
Rk256	XI2/XI0/XI1/net2#4	XI2/XI0/XI1/net2#5	31.000000
+ $metal1_conn
Rk257	XI2/XI0/XI1/net2#7	XI2/XI0/XI1/net2#8	31.000000
+ $metal1_conn
Rk258	XI2/XI1/D#17	XI2/XI1/D#2	0.292025	$metal1_conn
Rk259	XI2/XI1/D#2	XI2/XI1/D#19	0.466581	$metal1_conn
Rk260	net14#5	net14#17	45.731133	$metal1_conn
Rk261	SOUT2#11	SOUT2#8	0.156463	$metal1_conn
Rk262	SOUT2#8	SOUT2#2	45.836899	$metal1_conn
Rk263	VDD#69	VDD#70	15.500000	$metal1_conn
Rk264	GND#59	GND#60	37.500000	$metal1_conn
Rk265	VDD#71	VDD#72	31.001158	$metal1_conn
Rk266	XI2/XI1/XI4/net24#4	XI2/XI1/XI4/net24#2	45.402275
+ $metal1_conn
Rk267	XI2/XI1/XI4/net24#2	XI2/XI1/XI4/net24#9	0.668824
+ $metal1_conn
Rk268	XI2/XI1/D#20	XI2/XI1/D#4	45.082287	$metal1_conn
Rk269	XI2/XI1/XI4/net24#10	XI2/XI1/XI4/net24#11	15.500000
+ $metal1_conn
Rk270	XI2/XI1/XI4/net24#12	XI2/XI1/XI4/net24#13	0.688239
+ $metal1_conn
Rk271	XI2/XI1/Q#8	XI2/XI1/Q#9	37.500000	$metal1_conn
Rk272	XI2/XI0/XI1/net2#11	XI2/XI0/XI1/net2#12	0.001157
+ $metal1_conn
Rk273	XI2/XI0/XI1/net2#12	XI2/XI0/XI1/net2#13	0.169876
+ $metal1_conn
Rk274	XI2/XI0/XI1/net2#10	XI2/XI0/XI1/net2#11	37.500000
+ $metal1_conn
Rk275	XI2/net1#4	XI2/net1#2	46.295746	$metal1_conn
Rk276	XI2/XI0/XI0/BNOT#9	XI2/XI0/XI0/BNOT#10	2.761596
+ $metal1_conn
Rk277	XI2/XI0/XI0/BNOT#11	XI2/XI0/XI0/BNOT#2	45.782852
+ $metal1_conn
Rk279	XI2/net1#6	XI2/net1#9	0.322022	$metal1_conn
Rk280	XI2/net1#9	XI2/net1#11	0.257371	$metal1_conn
Rk282	XI2/net1#7	XI2/net1#6	15.500000	$metal1_conn
Rk283	XI2/net1#10	XI2/net1#11	15.500000	$metal1_conn
Rk285	XI2/net1#14	XI2/net1#16	0.305642	$metal1_conn
Rk286	XI2/net1#16	XI2/net1#18	0.240992	$metal1_conn
Rk288	XI2/net1#13	XI2/net1#14	37.500000	$metal1_conn
Rk289	XI2/net1#17	XI2/net1#18	37.500000	$metal1_conn
Rk290	net14#8	net14#19	46.508373	$metal1_conn
Rk291	net14#19	net14#20	0.688033	$metal1_conn
Rk292	net14#20	net14#21	1.364706	$metal1_conn
Rk293	VDD#73	VDD#74	31.000000	$metal1_conn
Rk294	VDD#75	VDD#76	31.000000	$metal1_conn
Rk295	GND#61	GND#62	75.000000	$metal1_conn
Rk296	GND#63	GND#64	75.000000	$metal1_conn
Rk297	XI2/XI1/Q#2	XI2/XI1/Q#11	45.453136	$metal1_conn
Rk298	XI2/XI1/Q#11	XI2/XI1/Q#12	0.376483	$metal1_conn
Rk299	XI2/XI0/XI1/net2#2	XI2/XI0/XI1/net2#15	45.440205
+ $metal1_conn
Rk300	XI2/XI0/XI1/net2#15	XI2/XI0/XI1/net2#16	0.343778
+ $metal1_conn
Rk301	XI2/XI0/XI0/BNOT#4	XI2/XI0/XI0/BNOT#14	45.156464
+ $metal1_conn
Rk302	SOUT2#14	SOUT2#15	31.001158	$metal1_conn
Rk303	VDD#77	VDD#78	15.500000	$metal1_conn
Rk304	GND#65	GND#66	37.500000	$metal1_conn
Rk305	net21#10	net21#11	31.001158	$metal1_conn
Rk306	SOUT2#16	SOUT2#17	75.001549	$metal1_conn
Rk307	net21#12	net21#13	75.001549	$metal1_conn
Rk308	SOUT2#18	SOUT2#19	1.205139	$metal1_conn
Rk309	SOUT2#20	SOUT2#5	46.880508	$metal1_conn
Rk310	SOUT2#22	SOUT2#10	0.248977	$metal1_conn
Rk311	SOUT2#10	SOUT2#24	0.776813	$metal1_conn
Rk312	net21#14	net21#15	0.885980	$metal1_conn
Rk313	VDD#79	VDD#80	31.000000	$metal1_conn
Rk314	GND#67	GND#68	75.000000	$metal1_conn
Rk315	XI3/XI1/D#5	XI3/XI1/D#6	37.501156	$metal1_conn
Rk316	VDD#81	VDD#82	31.000000	$metal1_conn
Rk317	VDD#83	VDD#84	31.001158	$metal1_conn
Rk318	GND#69	GND#70	75.000000	$metal1_conn
Rk319	XI3/XI0/XI0/ANOT#4	XI3/XI0/XI0/ANOT#5	31.001158
+ $metal1_conn
Rk320	XI3/XI0/XI0/ANOT#6	XI3/XI0/XI0/ANOT#7	75.001549
+ $metal1_conn
Rk321	XI3/XI1/XI4/PHINOT#4	XI3/XI1/XI4/PHINOT#5	31.001158
+ $metal1_conn
Rk322	XI3/XI1/XI4/PHINOT#6	XI3/XI1/XI4/PHINOT#7	75.001549
+ $metal1_conn
Rk323	VDD#85	VDD#86	31.000000	$metal1_conn
Rk324	XI3/XI1/XI5/net13#2	XI3/XI1/XI5/net13#3	0.001157
+ $metal1_conn
Rk325	XI3/XI1/XI5/net13#3	XI3/XI1/XI5/net13#5	0.232308
+ $metal1_conn
Rk327	XI3/XI1/XI5/net13	XI3/XI1/XI5/net13#2	37.500000
+ $metal1_conn
Rk328	XI3/XI1/XI5/net13#4	XI3/XI1/XI5/net13#5	37.500000
+ $metal1_conn
Rk329	GND#71	GND#72	75.000000	$metal1_conn
Rk330	XI3/XI1/D#7	XI3/XI1/D#9	0.001157	$metal1_conn
Rk331	XI3/XI1/D#9	XI3/XI1/D#10	0.120231	$metal1_conn
Rk332	XI3/XI1/D#10	XI3/XI1/D#12	0.114924	$metal1_conn
Rk334	XI3/XI1/D#8	XI3/XI1/D#9	31.000000	$metal1_conn
Rk335	XI3/XI1/D#11	XI3/XI1/D#12	31.000000	$metal1_conn
Rk336	XI3/XI0/XI0/BNOT#5	XI3/XI0/XI0/BNOT#6	31.001158
+ $metal1_conn
Rk337	GND#73	GND#74	37.500000	$metal1_conn
Rk338	VDD#87	VDD#88	31.000000	$metal1_conn
Rk339	XI3/XI0/XI0/BNOT#7	XI3/XI0/XI0/BNOT#8	75.001549
+ $metal1_conn
Rk340	XI3/XI1/D#14	XI3/XI1/D#15	0.450092	$metal1_conn
Rk341	XI3/XI1/D#15	XI3/XI1/D#16	0.266916	$metal1_conn
Rk342	GND#75	GND#76	37.500000	$metal1_conn
Rk343	VDD#89	VDD#90	31.000000	$metal1_conn
Rk344	XI3/XI1/Q#4	XI3/XI1/Q#5	15.500000	$metal1_conn
Rk345	XI3/XI1/XI4/net24#5	XI3/XI1/XI4/net24#6	37.500000
+ $metal1_conn
Rk346	XI3/XI1/XI4/PHINOT#2	XI3/XI1/XI4/PHINOT#9	46.516312
+ $metal1_conn
Rk347	VDD#91	VDD#92	15.500000	$metal1_conn
Rk348	GND#77	GND#78	37.500000	$metal1_conn
Rk349	VDD#93	VDD#94	15.500000	$metal1_conn
Rk350	GND#79	GND#80	37.500000	$metal1_conn
Rk351	XI3/XI1/Q#6	XI3/XI1/Q#7	0.365328	$metal1_conn
Rk352	XI3/XI0/XI0/ANOT#2	XI3/XI0/XI0/ANOT#9	46.855549
+ $metal1_conn
Rk354	XI3/XI0/XI1/XI0/net13#2	XI3/XI0/XI1/XI0/net13#4
+ 0.232308	$metal1_conn
Rk355	XI3/XI0/XI1/XI0/net13#4	XI3/XI0/XI1/XI0/net13#5
+ 37.501156	$metal1_conn
Rk356	XI3/XI0/XI1/XI0/net13	XI3/XI0/XI1/XI0/net13#2	37.500000
+ $metal1_conn
Rk358	XI3/XI0/XI1/net2#5	XI3/XI0/XI1/net2#8	0.237615
+ $metal1_conn
Rk359	XI3/XI0/XI1/net2#8	XI3/XI0/XI1/net2#9	0.001157
+ $metal1_conn
Rk360	XI3/XI0/XI1/net2#4	XI3/XI0/XI1/net2#5	31.000000
+ $metal1_conn
Rk361	XI3/XI0/XI1/net2#7	XI3/XI0/XI1/net2#8	31.000000
+ $metal1_conn
Rk362	XI3/XI1/D#17	XI3/XI1/D#2	0.292025	$metal1_conn
Rk363	XI3/XI1/D#2	XI3/XI1/D#19	0.466581	$metal1_conn
Rk364	net21#5	net21#17	45.731133	$metal1_conn
Rk365	SOUT3#11	SOUT3#8	0.156463	$metal1_conn
Rk366	SOUT3#8	SOUT3#2	45.836899	$metal1_conn
Rk367	VDD#95	VDD#96	15.500000	$metal1_conn
Rk368	GND#81	GND#82	37.500000	$metal1_conn
Rk369	VDD#97	VDD#98	31.001158	$metal1_conn
Rk370	XI3/XI1/XI4/net24#4	XI3/XI1/XI4/net24#2	45.402275
+ $metal1_conn
Rk371	XI3/XI1/XI4/net24#2	XI3/XI1/XI4/net24#9	0.668824
+ $metal1_conn
Rk372	XI3/XI1/D#20	XI3/XI1/D#4	45.082287	$metal1_conn
Rk373	XI3/XI1/XI4/net24#10	XI3/XI1/XI4/net24#11	15.500000
+ $metal1_conn
Rk374	XI3/XI1/XI4/net24#12	XI3/XI1/XI4/net24#13	0.688239
+ $metal1_conn
Rk375	XI3/XI1/Q#8	XI3/XI1/Q#9	37.500000	$metal1_conn
Rk376	XI3/XI0/XI1/net2#11	XI3/XI0/XI1/net2#12	0.001157
+ $metal1_conn
Rk377	XI3/XI0/XI1/net2#12	XI3/XI0/XI1/net2#13	0.169876
+ $metal1_conn
Rk378	XI3/XI0/XI1/net2#10	XI3/XI0/XI1/net2#11	37.500000
+ $metal1_conn
Rk379	XI3/net1#4	XI3/net1#2	46.295746	$metal1_conn
Rk380	XI3/XI0/XI0/BNOT#9	XI3/XI0/XI0/BNOT#10	2.761596
+ $metal1_conn
Rk381	XI3/XI0/XI0/BNOT#11	XI3/XI0/XI0/BNOT#2	45.782852
+ $metal1_conn
Rk383	XI3/net1#6	XI3/net1#9	0.322022	$metal1_conn
Rk384	XI3/net1#9	XI3/net1#11	0.257371	$metal1_conn
Rk386	XI3/net1#7	XI3/net1#6	15.500000	$metal1_conn
Rk387	XI3/net1#10	XI3/net1#11	15.500000	$metal1_conn
Rk389	XI3/net1#14	XI3/net1#16	0.305642	$metal1_conn
Rk390	XI3/net1#16	XI3/net1#18	0.240992	$metal1_conn
Rk392	XI3/net1#13	XI3/net1#14	37.500000	$metal1_conn
Rk393	XI3/net1#17	XI3/net1#18	37.500000	$metal1_conn
Rk394	net21#8	net21#19	46.508373	$metal1_conn
Rk395	net21#19	net21#20	0.688033	$metal1_conn
Rk396	net21#20	net21#21	1.364706	$metal1_conn
Rk397	VDD#99	VDD#100	31.000000	$metal1_conn
Rk398	VDD#101	VDD#102	31.000000	$metal1_conn
Rk399	GND#83	GND#84	75.000000	$metal1_conn
Rk400	GND#85	GND#86	75.000000	$metal1_conn
Rk401	XI3/XI1/Q#2	XI3/XI1/Q#11	45.453136	$metal1_conn
Rk402	XI3/XI1/Q#11	XI3/XI1/Q#12	0.376483	$metal1_conn
Rk403	XI3/XI0/XI1/net2#2	XI3/XI0/XI1/net2#15	45.440205
+ $metal1_conn
Rk404	XI3/XI0/XI1/net2#15	XI3/XI0/XI1/net2#16	0.343778
+ $metal1_conn
Rk405	XI3/XI0/XI0/BNOT#4	XI3/XI0/XI0/BNOT#14	45.156464
+ $metal1_conn
Rk406	SOUT3#14	SOUT3#15	31.001158	$metal1_conn
Rk407	VDD#103	VDD#104	15.500000	$metal1_conn
Rk408	GND#87	GND#88	37.500000	$metal1_conn
Rk409	COUT#1	COUT#2	31.001158	$metal1_conn
Rk410	SOUT3#16	SOUT3#17	75.001549	$metal1_conn
Rk411	COUT#3	COUT#4	75.001549	$metal1_conn
Rk412	SOUT3#18	SOUT3#19	1.205139	$metal1_conn
Rk413	SOUT3#20	SOUT3#5	46.880508	$metal1_conn
Rk414	SOUT3#22	SOUT3#10	0.248977	$metal1_conn
Rk415	SOUT3#10	SOUT3#24	0.776813	$metal1_conn
Rk416	COUT#5	COUT#6	0.885980	$metal1_conn
Rk417	VDD#105	VDD#107	0.045855	$metal1_conn
Rk418	VDD#107	VDD#108	0.256720	$metal1_conn
Rk419	VDD#108	VDD#109	0.194163	$metal1_conn
Rk420	VDD#109	VDD#110	0.085599	$metal1_conn
Rk421	VDD#110	VDD#111	0.390413	$metal1_conn
Rk422	VDD#111	VDD#112	0.275586	$metal1_conn
Rk423	VDD#112	VDD#114	0.045855	$metal1_conn
Rk424	VDD#114	VDD#115	0.256720	$metal1_conn
Rk425	VDD#115	VDD#116	0.194163	$metal1_conn
Rk426	VDD#116	VDD#117	0.085599	$metal1_conn
Rk427	VDD#117	VDD#118	0.390413	$metal1_conn
Rk428	VDD#118	VDD#119	0.275586	$metal1_conn
Rk429	VDD#119	VDD#121	0.045855	$metal1_conn
Rk430	VDD#121	VDD#122	0.256720	$metal1_conn
Rk431	VDD#122	VDD#123	0.194163	$metal1_conn
Rk432	VDD#123	VDD#124	0.085599	$metal1_conn
Rk433	VDD#124	VDD#125	0.390413	$metal1_conn
Rk434	VDD#125	VDD#126	0.275586	$metal1_conn
Rk435	VDD#126	VDD#128	0.045855	$metal1_conn
Rk436	VDD#128	VDD#129	0.256720	$metal1_conn
Rk437	VDD#129	VDD#130	0.194163	$metal1_conn
Rk438	VDD#130	VDD#131	0.085599	$metal1_conn
Rk439	VDD#131	VDD	0.315253	$metal1_conn
Rk440	VDD	VDD#132	0.075160	$metal1_conn
Rk441	VDD#106	VDD#107	18.750000	$metal1_conn
Rk442	VDD#113	VDD#114	18.750000	$metal1_conn
Rk443	VDD#120	VDD#121	18.750000	$metal1_conn
Rk444	VDD#127	VDD#128	18.750000	$metal1_conn
Rk445	VDD#133	VDD#135	0.047483	$metal1_conn
Rk446	VDD#135	VDD#136	0.214504	$metal1_conn
Rk447	VDD#136	VDD#137	0.041755	$metal1_conn
Rk448	VDD#137	VDD#138	0.185811	$metal1_conn
Rk449	VDD#138	VDD#139	0.085599	$metal1_conn
Rk450	VDD#139	VDD#140	0.081423	$metal1_conn
Rk451	VDD#140	VDD#141	0.151363	$metal1_conn
Rk452	VDD#141	VDD#142	0.044887	$metal1_conn
Rk453	VDD#142	VDD#143	0.125266	$metal1_conn
Rk454	VDD#143	VDD#144	0.273498	$metal1_conn
Rk455	VDD#144	VDD#146	0.047483	$metal1_conn
Rk456	VDD#146	VDD#147	0.214504	$metal1_conn
Rk457	VDD#147	VDD#148	0.041755	$metal1_conn
Rk458	VDD#148	VDD#149	0.185811	$metal1_conn
Rk459	VDD#149	VDD#150	0.085599	$metal1_conn
Rk460	VDD#150	VDD#151	0.081423	$metal1_conn
Rk461	VDD#151	VDD#152	0.151363	$metal1_conn
Rk462	VDD#152	VDD#153	0.044887	$metal1_conn
Rk463	VDD#153	VDD#154	0.125266	$metal1_conn
Rk464	VDD#154	VDD#155	0.273498	$metal1_conn
Rk465	VDD#155	VDD#157	0.047483	$metal1_conn
Rk466	VDD#157	VDD#158	0.214504	$metal1_conn
Rk467	VDD#158	VDD#159	0.041755	$metal1_conn
Rk468	VDD#159	VDD#160	0.185811	$metal1_conn
Rk469	VDD#160	VDD#161	0.085599	$metal1_conn
Rk470	VDD#161	VDD#162	0.081423	$metal1_conn
Rk471	VDD#162	VDD#163	0.151363	$metal1_conn
Rk472	VDD#163	VDD#164	0.044887	$metal1_conn
Rk473	VDD#164	VDD#165	0.125266	$metal1_conn
Rk474	VDD#165	VDD#166	0.273498	$metal1_conn
Rk475	VDD#166	VDD#168	0.047483	$metal1_conn
Rk476	VDD#168	VDD#169	0.214504	$metal1_conn
Rk477	VDD#169	VDD#170	0.041755	$metal1_conn
Rk478	VDD#170	VDD#171	0.185811	$metal1_conn
Rk479	VDD#171	VDD#172	0.085599	$metal1_conn
Rk480	VDD#172	VDD#173	0.081423	$metal1_conn
Rk481	VDD#173	VDD#174	0.151363	$metal1_conn
Rk482	VDD#174	VDD#175	0.044887	$metal1_conn
Rk483	VDD#175	VDD#176	0.625266	$metal1_conn
Rk484	VDD#134	VDD#135	18.750000	$metal1_conn
Rk485	VDD#145	VDD#146	18.750000	$metal1_conn
Rk486	VDD#156	VDD#157	18.750000	$metal1_conn
Rk487	VDD#167	VDD#168	18.750000	$metal1_conn
Rk488	GND#89	GND#91	0.156403	$metal1_conn
Rk489	GND#91	GND#92	0.045855	$metal1_conn
Rk490	GND#92	GND#93	0.167022	$metal1_conn
Rk491	GND#93	GND#94	0.313165	$metal1_conn
Rk492	GND#94	GND#95	0.277673	$metal1_conn
Rk493	GND#95	GND#96	0.129442	$metal1_conn
Rk494	GND#96	GND#98	0.315178	$metal1_conn
Rk495	GND#98	GND#99	0.045855	$metal1_conn
Rk496	GND#99	GND#100	0.167022	$metal1_conn
Rk497	GND#100	GND#101	0.313165	$metal1_conn
Rk498	GND#101	GND#102	0.277673	$metal1_conn
Rk499	GND#102	GND#103	0.129442	$metal1_conn
Rk500	GND#103	GND#105	0.315178	$metal1_conn
Rk501	GND#105	GND#106	0.045855	$metal1_conn
Rk502	GND#106	GND#107	0.167022	$metal1_conn
Rk503	GND#107	GND#108	0.313165	$metal1_conn
Rk504	GND#108	GND#109	0.277673	$metal1_conn
Rk505	GND#109	GND#110	0.129442	$metal1_conn
Rk506	GND#110	GND#112	0.315178	$metal1_conn
Rk507	GND#112	GND#113	0.045855	$metal1_conn
Rk508	GND#113	GND#114	0.167022	$metal1_conn
Rk509	GND#114	GND#115	0.313165	$metal1_conn
Rk510	GND#115	GND	0.200426	$metal1_conn
Rk511	GND	GND#116	0.077247	$metal1_conn
Rk512	GND#116	GND#117	0.129442	$metal1_conn
Rk513	GND#90	GND#91	15.500000	$metal1_conn
Rk514	GND#97	GND#98	15.500000	$metal1_conn
Rk515	GND#104	GND#105	15.500000	$metal1_conn
Rk516	GND#111	GND#112	15.500000	$metal1_conn
Rk517	COUT	COUT#7	0.367277	$metal1_conn
Rk518	PHI#25	PHI#26	1.759981	$metal1_conn
Rk519	PHI#26	PHI#27	1.695851	$metal1_conn
Rk520	PHI#27	PHI#28	2.331041	$metal1_conn
Rk521	PHI#28	PHI#29	1.695851	$metal1_conn
Rk522	PHI#29	PHI#30	2.331041	$metal1_conn
Rk523	PHI#30	PHI#31	1.695851	$metal1_conn
Rk524	PHI#31	PHI#32	2.331041	$metal1_conn
Rk525	PHI#32	PHI#33	1.695851	$metal1_conn
Rk526	PHI#33	PHI	0.279811	$metal1_conn
Rk527	RST#13	RST#14	3.362283	$metal1_conn
Rk528	RST#14	RST#15	3.932626	$metal1_conn
Rk529	RST#15	RST#16	3.932626	$metal1_conn
Rk530	RST#16	RST#17	3.932626	$metal1_conn
Rk531	RST#17	RST	0.214442	$metal1_conn
Rk532	GND#118	GND#119	15.548018	$metal1_conn
Rk533	GND#119	GND#120	0.210865	$metal1_conn
Rk534	GND#120	GND#121	0.194163	$metal1_conn
Rk535	GND#121	GND#122	0.085599	$metal1_conn
Rk536	GND#122	GND#123	0.070984	$metal1_conn
Rk537	GND#123	GND#124	0.151363	$metal1_conn
Rk538	GND#124	GND#125	0.168065	$metal1_conn
Rk539	GND#125	GND#127	0.323604	$metal1_conn
Rk540	GND#127	GND#128	0.048019	$metal1_conn
Rk541	GND#128	GND#129	0.210865	$metal1_conn
Rk542	GND#129	GND#130	0.194163	$metal1_conn
Rk543	GND#130	GND#131	0.085599	$metal1_conn
Rk544	GND#131	GND#132	0.070984	$metal1_conn
Rk545	GND#132	GND#133	0.151363	$metal1_conn
Rk546	GND#133	GND#134	0.168065	$metal1_conn
Rk547	GND#134	GND#136	0.323604	$metal1_conn
Rk548	GND#136	GND#137	0.048019	$metal1_conn
Rk549	GND#137	GND#138	0.210865	$metal1_conn
Rk550	GND#138	GND#139	0.194163	$metal1_conn
Rk551	GND#139	GND#140	0.085599	$metal1_conn
Rk552	GND#140	GND#141	0.070984	$metal1_conn
Rk553	GND#141	GND#142	0.151363	$metal1_conn
Rk554	GND#142	GND#143	0.168065	$metal1_conn
Rk555	GND#143	GND#145	0.323604	$metal1_conn
Rk556	GND#145	GND#146	0.048019	$metal1_conn
Rk557	GND#146	GND#147	0.210865	$metal1_conn
Rk558	GND#147	GND#148	0.194163	$metal1_conn
Rk559	GND#148	GND#149	0.085599	$metal1_conn
Rk560	GND#149	GND#150	0.070984	$metal1_conn
Rk561	GND#150	GND#151	0.151363	$metal1_conn
Rk562	GND#151	GND#152	0.168065	$metal1_conn
Rk563	GND#126	GND#127	15.500000	$metal1_conn
Rk564	GND#135	GND#136	15.500000	$metal1_conn
Rk565	GND#144	GND#145	15.500000	$metal1_conn
Rk596	net7#2	net7#20	45.000000	$metal1_conn
Rk614	net14#2	net14#20	45.000000	$metal1_conn
Rk632	net21#2	net21#20	45.000000	$metal1_conn
Rk638	PHI#23	PHI#26	45.000000	$metal1_conn
Rk639	PHI#20	PHI#27	45.000000	$metal1_conn
Rk640	PHI#17	PHI#28	45.000000	$metal1_conn
Rk641	PHI#14	PHI#29	45.000000	$metal1_conn
Rk642	PHI#11	PHI#30	45.000000	$metal1_conn
Rk643	PHI#8	PHI#31	45.000000	$metal1_conn
Rk644	PHI#5	PHI#32	45.000000	$metal1_conn
Rk645	PHI#2	PHI#33	45.000000	$metal1_conn
Rk646	RST#11	RST#14	45.000000	$metal1_conn
Rk647	RST#8	RST#15	45.000000	$metal1_conn
Rk648	RST#5	RST#16	45.000000	$metal1_conn
Rk649	RST#2	RST#17	45.000000	$metal1_conn
Rk577	CIN#2	CIN#12	45.000000	$metal1_conn
Rj1	GND#2	GND#117	1.222901	$metal2_conn
Rj2	XI0/XI1/D#6	XI0/XI1/D#16	1.047497	$metal2_conn
Rj3	VDD#132	VDD#4	0.992284	$metal2_conn
Rj4	GND#4	GND#152	1.208364	$metal2_conn
Rj5	VDD#2	VDD#176	0.479930	$metal2_conn
Rj6	VDD#176	VDD#5	0.463390	$metal2_conn
Rj7	XI0/XI0/XI0/ANOT#4	XI0/XI0/XI0/ANOT#9	0.904167
+ $metal2_conn
Rj8	XI0/XI0/XI0/ANOT#9	XI0/XI0/XI0/ANOT#6	0.844043
+ $metal2_conn
Rj9	XI0/XI1/XI4/PHINOT#4	XI0/XI1/XI4/PHINOT#9	0.676420
+ $metal2_conn
Rj10	XI0/XI1/XI4/PHINOT#9	XI0/XI1/XI4/PHINOT#6	1.071790
+ $metal2_conn
Rj11	XI0/XI1/D#15	XI0/XI1/D#10	1.725450	$metal2_conn
Rj12	VDD#175	VDD#8	0.982593	$metal2_conn
Rj13	GND#6	GND#116	1.222901	$metal2_conn
Rj14	XI0/XI0/XI0/BNOT#5	XI0/XI0/XI0/BNOT#10	0.812099
+ $metal2_conn
Rj15	XI0/XI0/XI0/BNOT#10	XI0/XI0/XI0/BNOT#7	0.936111
+ $metal2_conn
Rj16	GND#151	GND#8	0.968056	$metal2_conn
Rj17	VDD#10	VDD#174	0.969733	$metal2_conn
Rj18	XI0/XI1/D#19	XI0/XI1/D#14	1.901297	$metal2_conn
Rj19	CIN#11	CIN#13	2.327717	$metal2_conn
Rj20	GND#150	GND#10	0.968056	$metal2_conn
Rj21	VDD#12	VDD#173	0.969733	$metal2_conn
Rj22	XI0/XI1/Q#5	XI0/XI1/Q#7	0.828519	$metal2_conn
Rj23	XI0/XI1/XI4/net24#13	XI0/XI1/XI4/net24#9	0.691678
+ $metal2_conn
Rj24	XI0/XI1/XI4/net24#9	XI0/XI1/XI4/net24#6	0.509517
+ $metal2_conn
Rj25	VDD#131	VDD#14	0.901204	$metal2_conn
Rj26	GND#12	GND#149	0.968056	$metal2_conn
Rj27	VDD#172	VDD#16	0.906050	$metal2_conn
Rj28	GND#14	GND#115	0.972901	$metal2_conn
Rj29	XI0/XI1/Q#6	XI0/XI1/Q#12	1.452264	$metal2_conn
Rj30	XI0/XI0/XI1/net2#16	XI0/XI0/XI1/net2#5	1.013344
+ $metal2_conn
Rj31	XI0/XI1/D#20	XI0/XI1/D#17	1.635054	$metal2_conn
Rj32	SOUT0#11	SOUT0#24	1.576636	$metal2_conn
Rj33	VDD#130	VDD#18	0.901204	$metal2_conn
Rj34	GND#16	GND#148	0.968056	$metal2_conn
Rj35	VDD#20	VDD#171	0.969733	$metal2_conn
Rj36	XI0/XI1/XI4/net24#11	XI0/XI1/XI4/net24#12	1.124105
+ $metal2_conn
Rj37	XI0/XI1/Q#11	XI0/XI1/Q#9	1.098889	$metal2_conn
Rj38	XI0/XI0/XI1/net2#13	XI0/XI0/XI1/net2#15	1.755926
+ $metal2_conn
Rj39	XI0/net1#4	XI0/net1#23	1.154167	$metal2_conn
Rj40	XI0/net1#23	XI0/net1#16	1.449754	$metal2_conn
Rj41	XI0/XI0/XI0/BNOT#14	XI0/XI0/XI0/BNOT#9	0.800432
+ $metal2_conn
Rj42	XI0/XI0/XI0/BNOT#9	XI0/XI0/XI0/BNOT#11	0.679290
+ $metal2_conn
Rj43	VDD#129	VDD#22	0.992284	$metal2_conn
Rj44	GND#20	GND#170	0.725399	$metal2_conn
Rj45	GND#170	GND#18	0.703519	$metal2_conn
Rj46	VDD#24	VDD#170	0.988246	$metal2_conn
Rj47	SOUT0#14	SOUT0#19	1.112531	$metal2_conn
Rj48	SOUT0#19	SOUT0#16	0.635679	$metal2_conn
Rj49	VDD#169	VDD#26	0.906857	$metal2_conn
Rj50	GND#22	GND#114	0.972901	$metal2_conn
Rj51	net7#12	net7#15	0.756821	$metal2_conn
Rj52	net7#15	net7#10	0.991389	$metal2_conn
Rj53	SOUT0	SOUT0#18	1.201729	$metal2_conn
Rj54	SOUT0#18	SOUT0#20	0.919002	$metal2_conn
Rj55	SOUT0#20	SOUT0#22	2.494246	$metal2_conn
Rj56	net7#14	net7#21	2.719596	$metal2_conn
Rj57	GND#146	GND#113	3.873489	$metal2_conn
Rj58	VDD#126	VDD#166	3.912255	$metal2_conn
Rj59	GND#24	GND#110	1.222901	$metal2_conn
Rj60	XI1/XI1/D#6	XI1/XI1/D#16	1.047497	$metal2_conn
Rj61	VDD#125	VDD#30	0.992284	$metal2_conn
Rj62	GND#26	GND#143	1.208364	$metal2_conn
Rj63	VDD#28	VDD#207	0.479930	$metal2_conn
Rj64	VDD#207	VDD#31	0.463390	$metal2_conn
Rj65	XI1/XI0/XI0/ANOT#4	XI1/XI0/XI0/ANOT#9	0.904167
+ $metal2_conn
Rj66	XI1/XI0/XI0/ANOT#9	XI1/XI0/XI0/ANOT#6	0.844043
+ $metal2_conn
Rj67	XI1/XI1/XI4/PHINOT#4	XI1/XI1/XI4/PHINOT#9	0.676420
+ $metal2_conn
Rj68	XI1/XI1/XI4/PHINOT#9	XI1/XI1/XI4/PHINOT#6	1.071790
+ $metal2_conn
Rj69	XI1/XI1/D#15	XI1/XI1/D#10	1.725450	$metal2_conn
Rj70	VDD#164	VDD#34	0.982593	$metal2_conn
Rj71	GND#28	GND#109	1.222901	$metal2_conn
Rj72	XI1/XI0/XI0/BNOT#5	XI1/XI0/XI0/BNOT#10	0.812099
+ $metal2_conn
Rj73	XI1/XI0/XI0/BNOT#10	XI1/XI0/XI0/BNOT#7	0.936111
+ $metal2_conn
Rj74	GND#142	GND#30	0.968056	$metal2_conn
Rj75	VDD#36	VDD#163	0.969733	$metal2_conn
Rj76	XI1/XI1/D#19	XI1/XI1/D#14	1.901297	$metal2_conn
Rj77	net7#17	net7#19	2.327717	$metal2_conn
Rj78	GND#141	GND#32	0.968056	$metal2_conn
Rj79	VDD#38	VDD#162	0.969733	$metal2_conn
Rj80	XI1/XI1/Q#5	XI1/XI1/Q#7	0.828519	$metal2_conn
Rj81	XI1/XI1/XI4/net24#13	XI1/XI1/XI4/net24#9	0.691678
+ $metal2_conn
Rj82	XI1/XI1/XI4/net24#9	XI1/XI1/XI4/net24#6	0.509517
+ $metal2_conn
Rj83	VDD#124	VDD#40	0.901204	$metal2_conn
Rj84	GND#34	GND#140	0.968056	$metal2_conn
Rj85	VDD#161	VDD#42	0.906050	$metal2_conn
Rj86	GND#36	GND#108	0.972901	$metal2_conn
Rj87	XI1/XI1/Q#6	XI1/XI1/Q#12	1.452264	$metal2_conn
Rj88	XI1/XI0/XI1/net2#16	XI1/XI0/XI1/net2#5	1.013344
+ $metal2_conn
Rj89	XI1/XI1/D#20	XI1/XI1/D#17	1.635054	$metal2_conn
Rj90	SOUT1#11	SOUT1#24	1.576636	$metal2_conn
Rj91	VDD#123	VDD#44	0.901204	$metal2_conn
Rj92	GND#38	GND#139	0.968056	$metal2_conn
Rj93	VDD#46	VDD#160	0.969733	$metal2_conn
Rj94	XI1/XI1/XI4/net24#11	XI1/XI1/XI4/net24#12	1.124105
+ $metal2_conn
Rj95	XI1/XI1/Q#11	XI1/XI1/Q#9	1.098889	$metal2_conn
Rj96	XI1/XI0/XI1/net2#13	XI1/XI0/XI1/net2#15	1.755926
+ $metal2_conn
Rj97	XI1/net1#4	XI1/net1#23	1.154167	$metal2_conn
Rj98	XI1/net1#23	XI1/net1#16	1.449754	$metal2_conn
Rj99	XI1/XI0/XI0/BNOT#14	XI1/XI0/XI0/BNOT#9	0.800432
+ $metal2_conn
Rj100	XI1/XI0/XI0/BNOT#9	XI1/XI0/XI0/BNOT#11	0.679290
+ $metal2_conn
Rj101	VDD#122	VDD#48	0.992284	$metal2_conn
Rj102	GND#42	GND#193	0.725399	$metal2_conn
Rj103	GND#193	GND#40	0.703519	$metal2_conn
Rj104	VDD#50	VDD#159	0.988246	$metal2_conn
Rj105	SOUT1#14	SOUT1#19	1.112531	$metal2_conn
Rj106	SOUT1#19	SOUT1#16	0.635679	$metal2_conn
Rj107	VDD#158	VDD#52	0.906857	$metal2_conn
Rj108	GND#44	GND#107	0.972901	$metal2_conn
Rj109	net14#12	net14#15	0.756821	$metal2_conn
Rj110	net14#15	net14#10	0.991389	$metal2_conn
Rj111	SOUT1	SOUT1#18	1.201729	$metal2_conn
Rj112	SOUT1#18	SOUT1#20	0.919002	$metal2_conn
Rj113	SOUT1#20	SOUT1#22	2.494246	$metal2_conn
Rj114	net14#14	net14#21	2.719596	$metal2_conn
Rj115	GND#137	GND#106	3.873489	$metal2_conn
Rj116	VDD#119	VDD#155	3.912255	$metal2_conn
Rj117	GND#46	GND#103	1.222901	$metal2_conn
Rj118	XI2/XI1/D#6	XI2/XI1/D#16	1.047497	$metal2_conn
Rj119	VDD#118	VDD#56	0.992284	$metal2_conn
Rj120	GND#48	GND#134	1.208364	$metal2_conn
Rj121	VDD#54	VDD#234	0.479930	$metal2_conn
Rj122	VDD#234	VDD#57	0.463390	$metal2_conn
Rj123	XI2/XI0/XI0/ANOT#4	XI2/XI0/XI0/ANOT#9	0.904167
+ $metal2_conn
Rj124	XI2/XI0/XI0/ANOT#9	XI2/XI0/XI0/ANOT#6	0.844043
+ $metal2_conn
Rj125	XI2/XI1/XI4/PHINOT#4	XI2/XI1/XI4/PHINOT#9	0.676420
+ $metal2_conn
Rj126	XI2/XI1/XI4/PHINOT#9	XI2/XI1/XI4/PHINOT#6	1.071790
+ $metal2_conn
Rj127	XI2/XI1/D#15	XI2/XI1/D#10	1.725450	$metal2_conn
Rj128	VDD#153	VDD#60	0.982593	$metal2_conn
Rj129	GND#50	GND#102	1.222901	$metal2_conn
Rj130	XI2/XI0/XI0/BNOT#5	XI2/XI0/XI0/BNOT#10	0.812099
+ $metal2_conn
Rj131	XI2/XI0/XI0/BNOT#10	XI2/XI0/XI0/BNOT#7	0.936111
+ $metal2_conn
Rj132	GND#133	GND#52	0.968056	$metal2_conn
Rj133	VDD#62	VDD#152	0.969733	$metal2_conn
Rj134	XI2/XI1/D#19	XI2/XI1/D#14	1.901297	$metal2_conn
Rj135	net14#17	net14#19	2.327717	$metal2_conn
Rj136	GND#132	GND#54	0.968056	$metal2_conn
Rj137	VDD#64	VDD#151	0.969733	$metal2_conn
Rj138	XI2/XI1/Q#5	XI2/XI1/Q#7	0.828519	$metal2_conn
Rj139	XI2/XI1/XI4/net24#13	XI2/XI1/XI4/net24#9	0.691678
+ $metal2_conn
Rj140	XI2/XI1/XI4/net24#9	XI2/XI1/XI4/net24#6	0.509517
+ $metal2_conn
Rj141	VDD#117	VDD#66	0.901204	$metal2_conn
Rj142	GND#56	GND#131	0.968056	$metal2_conn
Rj143	VDD#150	VDD#68	0.906050	$metal2_conn
Rj144	GND#58	GND#101	0.972901	$metal2_conn
Rj145	XI2/XI1/Q#6	XI2/XI1/Q#12	1.452264	$metal2_conn
Rj146	XI2/XI0/XI1/net2#16	XI2/XI0/XI1/net2#5	1.013344
+ $metal2_conn
Rj147	XI2/XI1/D#20	XI2/XI1/D#17	1.635054	$metal2_conn
Rj148	SOUT2#11	SOUT2#24	1.576636	$metal2_conn
Rj149	VDD#116	VDD#70	0.901204	$metal2_conn
Rj150	GND#60	GND#130	0.968056	$metal2_conn
Rj151	VDD#72	VDD#149	0.969733	$metal2_conn
Rj152	XI2/XI1/XI4/net24#11	XI2/XI1/XI4/net24#12	1.124105
+ $metal2_conn
Rj153	XI2/XI1/Q#11	XI2/XI1/Q#9	1.098889	$metal2_conn
Rj154	XI2/XI0/XI1/net2#13	XI2/XI0/XI1/net2#15	1.755926
+ $metal2_conn
Rj155	XI2/net1#4	XI2/net1#23	1.154167	$metal2_conn
Rj156	XI2/net1#23	XI2/net1#16	1.449754	$metal2_conn
Rj157	XI2/XI0/XI0/BNOT#14	XI2/XI0/XI0/BNOT#9	0.800432
+ $metal2_conn
Rj158	XI2/XI0/XI0/BNOT#9	XI2/XI0/XI0/BNOT#11	0.679290
+ $metal2_conn
Rj159	VDD#115	VDD#74	0.992284	$metal2_conn
Rj160	GND#64	GND#216	0.725399	$metal2_conn
Rj161	GND#216	GND#62	0.703519	$metal2_conn
Rj162	VDD#76	VDD#148	0.988246	$metal2_conn
Rj163	SOUT2#14	SOUT2#19	1.112531	$metal2_conn
Rj164	SOUT2#19	SOUT2#16	0.635679	$metal2_conn
Rj165	VDD#147	VDD#78	0.906857	$metal2_conn
Rj166	GND#66	GND#100	0.972901	$metal2_conn
Rj167	net21#12	net21#15	0.756821	$metal2_conn
Rj168	net21#15	net21#10	0.991389	$metal2_conn
Rj169	SOUT2	SOUT2#18	1.201729	$metal2_conn
Rj170	SOUT2#18	SOUT2#20	0.919002	$metal2_conn
Rj171	SOUT2#20	SOUT2#22	2.494246	$metal2_conn
Rj172	net21#14	net21#21	2.719596	$metal2_conn
Rj173	GND#128	GND#99	3.873489	$metal2_conn
Rj174	VDD#112	VDD#144	3.912255	$metal2_conn
Rj175	GND#68	GND#96	1.222901	$metal2_conn
Rj176	XI3/XI1/D#6	XI3/XI1/D#16	1.047497	$metal2_conn
Rj177	VDD#111	VDD#82	0.992284	$metal2_conn
Rj178	GND#70	GND#125	1.208364	$metal2_conn
Rj179	VDD#80	VDD#261	0.479930	$metal2_conn
Rj180	VDD#261	VDD#83	0.463390	$metal2_conn
Rj181	XI3/XI0/XI0/ANOT#4	XI3/XI0/XI0/ANOT#9	0.904167
+ $metal2_conn
Rj182	XI3/XI0/XI0/ANOT#9	XI3/XI0/XI0/ANOT#6	0.844043
+ $metal2_conn
Rj183	XI3/XI1/XI4/PHINOT#4	XI3/XI1/XI4/PHINOT#9	0.676420
+ $metal2_conn
Rj184	XI3/XI1/XI4/PHINOT#9	XI3/XI1/XI4/PHINOT#6	1.071790
+ $metal2_conn
Rj185	XI3/XI1/D#15	XI3/XI1/D#10	1.725450	$metal2_conn
Rj186	VDD#142	VDD#86	0.982593	$metal2_conn
Rj187	GND#72	GND#95	1.222901	$metal2_conn
Rj188	XI3/XI0/XI0/BNOT#5	XI3/XI0/XI0/BNOT#10	0.812099
+ $metal2_conn
Rj189	XI3/XI0/XI0/BNOT#10	XI3/XI0/XI0/BNOT#7	0.936111
+ $metal2_conn
Rj190	GND#124	GND#74	0.968056	$metal2_conn
Rj191	VDD#88	VDD#141	0.969733	$metal2_conn
Rj192	XI3/XI1/D#19	XI3/XI1/D#14	1.901297	$metal2_conn
Rj193	net21#17	net21#19	2.327717	$metal2_conn
Rj194	GND#123	GND#76	0.968056	$metal2_conn
Rj195	VDD#90	VDD#140	0.969733	$metal2_conn
Rj196	XI3/XI1/Q#5	XI3/XI1/Q#7	0.828519	$metal2_conn
Rj197	XI3/XI1/XI4/net24#13	XI3/XI1/XI4/net24#9	0.691678
+ $metal2_conn
Rj198	XI3/XI1/XI4/net24#9	XI3/XI1/XI4/net24#6	0.509517
+ $metal2_conn
Rj199	VDD#110	VDD#92	0.901204	$metal2_conn
Rj200	GND#78	GND#122	0.968056	$metal2_conn
Rj201	VDD#139	VDD#94	0.906050	$metal2_conn
Rj202	GND#80	GND#94	0.972901	$metal2_conn
Rj203	XI3/XI1/Q#6	XI3/XI1/Q#12	1.452264	$metal2_conn
Rj204	XI3/XI0/XI1/net2#16	XI3/XI0/XI1/net2#5	1.013344
+ $metal2_conn
Rj205	XI3/XI1/D#20	XI3/XI1/D#17	1.635054	$metal2_conn
Rj206	SOUT3#11	SOUT3#24	1.576636	$metal2_conn
Rj207	VDD#109	VDD#96	0.901204	$metal2_conn
Rj208	GND#82	GND#121	0.968056	$metal2_conn
Rj209	VDD#98	VDD#138	0.969733	$metal2_conn
Rj210	XI3/XI1/XI4/net24#11	XI3/XI1/XI4/net24#12	1.124105
+ $metal2_conn
Rj211	XI3/XI1/Q#11	XI3/XI1/Q#9	1.098889	$metal2_conn
Rj212	XI3/XI0/XI1/net2#13	XI3/XI0/XI1/net2#15	1.755926
+ $metal2_conn
Rj213	XI3/net1#4	XI3/net1#23	1.154167	$metal2_conn
Rj214	XI3/net1#23	XI3/net1#16	1.449754	$metal2_conn
Rj215	XI3/XI0/XI0/BNOT#14	XI3/XI0/XI0/BNOT#9	0.800432
+ $metal2_conn
Rj216	XI3/XI0/XI0/BNOT#9	XI3/XI0/XI0/BNOT#11	0.679290
+ $metal2_conn
Rj217	VDD#108	VDD#100	0.992284	$metal2_conn
Rj218	GND#86	GND#239	0.725399	$metal2_conn
Rj219	GND#239	GND#84	0.703519	$metal2_conn
Rj220	VDD#102	VDD#137	0.988246	$metal2_conn
Rj221	SOUT3#14	SOUT3#19	1.112531	$metal2_conn
Rj222	SOUT3#19	SOUT3#16	0.635679	$metal2_conn
Rj223	VDD#136	VDD#104	0.906857	$metal2_conn
Rj224	GND#88	GND#93	0.972901	$metal2_conn
Rj225	COUT#3	COUT#6	0.756821	$metal2_conn
Rj226	COUT#6	COUT#1	0.991389	$metal2_conn
Rj227	SOUT3	SOUT3#18	1.201729	$metal2_conn
Rj228	SOUT3#18	SOUT3#20	0.919002	$metal2_conn
Rj229	SOUT3#20	SOUT3#22	2.494246	$metal2_conn
Rj230	COUT#5	COUT#7	2.719596	$metal2_conn
Rj231	GND#119	GND#92	3.873489	$metal2_conn
Rj232	VDD#105	VDD#133	3.912255	$metal2_conn
Rj315	XI0/net1#9	XI0/net1#23	0.500000	$metal2_conn
Rj587	VDD#143	VDD#261	0.500000	$metal2_conn
Rj325	GND#147	GND#170	0.500000	$metal2_conn
Rj472	VDD#154	VDD#234	0.500000	$metal2_conn
Rj357	VDD#165	VDD#207	0.500000	$metal2_conn
Rj660	XI3/net1#9	XI3/net1#23	0.500000	$metal2_conn
Rj670	GND#120	GND#239	0.500000	$metal2_conn
Rj545	XI2/net1#9	XI2/net1#23	0.500000	$metal2_conn
Rj555	GND#129	GND#216	0.500000	$metal2_conn
Rj430	XI1/net1#9	XI1/net1#23	0.500000	$metal2_conn
Rj440	GND#138	GND#193	0.500000	$metal2_conn
*
*       CAPACITOR CARDS
*
*
C1	SOUT2#18	PHI#17	1.77809e-17
C2	GND#120	SOUT3#16	1.37047e-17
C3	XI3/XI1/Q#5	XI3/XI1/Q#4	9.30041e-18
C4	XI3/XI1/XI4/PHINOT#6	XI3/XI1/XI4/PHINOT#7	4.46757e-18
C5	GND#14	XI0/XI0/XI0/ANOT#3	2.55369e-18
C6	VDD#150	XI2/XI0/XI0/ANOT	1.82797e-18
C7	net21#19	SOUT3#8	2.94542e-17
C8	GND#147	SOUT0#16	1.37047e-17
C9	XI0/XI1/XI4/net24#13	XI0/XI1/Q#7	3.21387e-18
C10	GND#28	SOUT1#3	4.36955e-18
C11	VDD#124	XI1/XI1/XI4/net24	4.3074e-18
C12	XI0/XI1/Q#5	XI0/XI1/XI4/PHINOT	8.79316e-18
C13	GND#107	net7#9	4.17672e-18
C14	XI1/XI1/XI4/net24	XI1/XI1/D#3	2.28624e-18
C15	XI0/XI1/D#20	XI0/XI1/XI4/net24#11	1.30924e-17
C16	XI3/XI1/Q#6	VDD#109	1.9494e-18
C17	RST#13	GND#118	1.50587e-17
C18	PHI#12	XI1/XI1/Q#3	3.05252e-18
C19	GND#128	VDD#145	1.10177e-17
C20	SOUT1#16	SOUT1#18	1.30402e-17
C21	VDD#16	XI0/net1#9	2.69821e-18
C22	VDD#175	VDD	1.8633e-17
C23	VDD#164	VDD#163	1.68962e-17
C24	VDD#110	VDD	8.4118e-17
C25	XI3/XI0/XI0/BNOT#11	net21#9	3.59305e-18
C26	net14#21	VDD#158	6.72863e-18
C27	SOUT3#18	XI3/XI1/Q#3	1.55626e-18
C28	XI0/XI1/XI4/net24#9	XI0/XI1/XI4/PHINOT#2	1.74823e-18
C29	XI3/XI1/Q#6	XI3/XI1/XI4/PHINOT#2	2.75539e-18
C30	XI0/XI0/XI0/ANOT	CIN#7	1.29274e-18
C31	COUT#6	XI3/XI0/XI1/net2	7.48119e-18
C32	net21#10	XI2/XI0/XI1/net2#2	5.88268e-18
C33	net21#10	XI2/XI0/XI1/net2#3	6.65581e-18
C34	GND#58	XI2/XI0/XI0/BNOT#2	1.48416e-18
C35	GND#113	net7#21	1.0327e-16
C36	SOUT1#8	VDD#42	1.33308e-17
C37	XI0/XI1/Q#11	PHI#5	1.16343e-17
C38	net14#19	XI2/XI0/XI0/ANOT#2	1.52499e-17
C39	SOUT0#18	GND#146	3.44305e-17
C40	GND#151	XI0/net1	4.15538e-18
C41	GND#44	GND#106	8.15798e-18
C42	XI1/net1#16	XI1/XI0/XI0/BNOT#9	1.54391e-17
C43	SOUT0#11	XI0/net1#9	2.44574e-17
C44	XI1/XI1/XI4/net24#13	PHI#11	9.76906e-18
C45	XI0/XI0/XI1/net2#16	XI0/net1#4	3.40431e-17
C46	XI0/XI1/Q#11	XI0/XI1/XI4/net24#12	2.96161e-17
C47	XI1/XI0/XI0/ANOT#2	net7#8	2.9337e-18
C48	GND#88	GND#87	7.74457e-18
C49	VDD#136	COUT#1	1.49363e-17
C50	VDD#139	VDD	1.44935e-17
C51	GND#132	XI2/XI1/XI4/PHINOT#3	3.59673e-18
C52	VDD#26	CIN#7	4.04071e-18
C53	XI0/XI0/XI0/BNOT#5	VDD	8.81368e-18
C54	XI0/net1#2	SOUT0#6	1.96305e-17
C55	XI2/XI1/Q#5	VDD#66	6.36626e-17
C56	XI1/XI1/D#10	net7#17	1.25206e-17
C57	VDD#74	SOUT2	4.09262e-18
C58	XI0/net1#4	VDD#171	1.4412e-17
C59	SOUT3#22	COUT#7	1.19768e-16
C60	XI2/XI1/Q#7	VDD#117	1.95651e-18
C61	PHI#22	XI3/XI1/Q	2.93097e-18
C62	GND#93	SOUT3#22	9.0763e-18
C63	VDD#174	VDD	1.94359e-17
C64	SOUT2	VDD#115	3.80499e-17
C65	GND#129	XI2/XI1/Q#3	2.16945e-18
C66	XI3/XI1/Q#6	VDD	9.99629e-18
C67	net21#6	XI3/XI0/XI1/net2#3	1.19235e-18
C68	VDD#174	VDD#10	1.0238e-17
C69	VDD#144	RST#11	2.35653e-17
C70	XI2/XI1/D#6	XI2/XI1/D#5	4.49187e-18
C71	GND#86	SOUT3#20	5.19922e-18
C72	XI2/XI1/XI4/net24#9	XI2/XI1/D#2	3.0624e-17
C73	XI2/XI0/XI0/BNOT#7	SOUT2#3	5.63912e-18
C74	net21#17	VDD#90	1.45914e-17
C75	SOUT1#24	XI1/XI0/XI0/ANOT#3	2.93467e-18
C76	XI2/net1#4	net14#5	1.24619e-17
C77	VDD#151	SOUT2#6	4.21273e-18
C78	net7#17	VDD#38	1.45914e-17
C79	VDD#96	VDD#109	1.16687e-17
C80	XI0/net1#9	XI0/XI0/XI0/BNOT#9	3.86468e-18
C81	CIN#13	VDD#16	1.37441e-17
C82	XI2/XI1/D#16	XI2/XI1/D#15	9.36359e-18
C83	XI3/XI1/XI4/net24#13	PHI#23	9.76906e-18
C84	net14#19	VDD#152	1.34565e-17
C85	VDD#126	XI0/XI1/Q#2	2.47832e-18
C86	XI1/XI1/D#10	RST#6	3.88703e-18
C87	XI3/XI0/XI1/net2#16	VDD	3.04753e-18
C88	XI3/XI0/XI1/net2#15	SOUT3#20	5.36179e-18
C89	XI1/XI0/XI0/ANOT#4	XI1/XI0/XI0/BNOT#10	2.24348e-18
C90	XI2/XI0/XI0/BNOT#7	XI2/XI0/XI0/BNOT#8	4.0203e-18
C91	XI2/XI1/XI4/net24#13	XI2/XI1/XI4/PHINOT#2	2.64065e-17
C92	XI0/XI0/XI1/net2#15	SOUT0#20	5.36179e-18
C93	XI3/XI1/XI4/net24#12	XI3/XI1/Q#2	2.89847e-18
C94	RST#11	GND#74	1.03647e-17
C95	XI2/XI1/D#20	XI2/XI1/XI4/net24#12	1.97297e-17
C96	XI3/XI1/XI4/PHINOT#4	XI3/XI1/XI4/PHINOT#5	5.34824e-18
C97	CIN#13	VDD	7.38122e-18
C98	net14#19	SOUT2#2	6.17276e-17
C99	XI1/net1#4	net7#5	1.24619e-17
C100	XI0/XI1/D#15	XI0/net1#2	3.59645e-18
C101	XI1/XI1/Q#12	XI1/XI1/XI4/net24#13	1.81832e-17
C102	CIN#11	VDD	6.33291e-18
C103	GND#119	XI3/XI0/XI1/net2#2	1.86055e-18
C104	XI1/XI0/XI0/ANOT#9	SOUT1#2	2.69483e-18
C105	XI3/XI0/XI1/net2#16	SOUT3#5	2.87586e-18
C106	XI3/XI1/D#20	VDD	3.67809e-18
C107	VDD#18	XI0/XI1/XI4/net24	1.58831e-18
C108	SOUT0#11	XI0/XI0/XI0/BNOT#14	3.25292e-18
C109	SOUT1#19	XI1/XI1/Q#2	6.59904e-18
C110	GND#117	GND#2	8.47392e-18
C111	GND#103	GND#46	8.47392e-18
C112	XI2/XI0/XI1/net2#15	net21#10	6.82353e-18
C113	XI0/XI1/Q#9	GND#18	1.37107e-17
C114	XI1/XI0/XI0/ANOT#9	net7#3	1.29853e-18
C115	XI3/XI1/D#20	XI3/XI1/XI4/net24#11	1.30924e-17
C116	XI2/XI1/XI4/net24#11	VDD#116	1.56401e-17
C117	VDD#158	XI1/XI0/XI1/net2#2	1.54384e-18
C118	XI3/XI0/XI1/net2#13	RST#11	2.21589e-17
C119	VDD#38	XI1/net1#2	1.29263e-17
C120	XI0/XI1/D#3	PHI#4	5.34502e-17
C121	XI3/XI0/XI0/ANOT#4	SOUT3#1	1.96312e-18
C122	VDD#173	VDD	2.56909e-17
C123	XI3/XI1/Q#11	XI3/XI1/XI4/net24#12	2.96161e-17
C124	SOUT2#14	SOUT2	3.64962e-17
C125	XI3/net1#9	XI3/XI0/XI0/BNOT#9	3.86468e-18
C126	XI3/XI0/XI0/BNOT#5	SOUT3#2	1.8238e-17
C127	GND#44	SOUT1#10	1.12163e-17
C128	GND#80	XI3/XI0/XI0/BNOT#2	1.48416e-18
C129	GND#102	XI2/XI0/XI0/BNOT#7	1.31853e-17
C130	GND#146	XI0/XI0/XI1/net2#2	1.86055e-18
C131	PHI#23	XI3/XI1/Q	1.18127e-17
C132	VDD#102	XI3/XI0/XI1/net2#2	8.46721e-18
C133	COUT#3	XI3/XI0/XI1/net2	5.18165e-18
C134	GND#94	GND#80	9.66245e-18
C135	XI3/net1#4	VDD#138	1.4412e-17
C136	SOUT2#11	XI2/XI0/XI0/ANOT#2	1.22267e-18
C137	VDD#78	SOUT2#22	3.78854e-17
C138	RST#12	XI3/net1#2	1.10422e-17
C139	XI3/XI0/XI0/ANOT#9	SOUT3#2	2.69483e-18
C140	XI1/XI1/D#2	XI1/XI1/D#17	3.60142e-18
C141	SOUT2#4	net14#4	4.68557e-18
C142	RST#2	GND#150	9.1293e-18
C143	VDD#14	XI0/XI1/D#3	1.58831e-18
C144	XI3/XI0/XI1/net2#16	XI3/net1#4	3.40431e-17
C145	VDD#64	SOUT2#6	4.07255e-18
C146	XI2/XI1/Q#11	PHI#17	1.16343e-17
C147	XI2/XI1/D#15	XI2/XI1/D#14	4.56509e-18
C148	XI0/XI1/Q#11	SOUT0#19	7.03151e-18
C149	XI1/XI1/D#15	XI1/net1	1.96101e-17
C150	XI3/XI1/XI4/PHINOT#6	XI3/XI1/D#19	8.37816e-18
C151	XI2/XI0/XI0/BNOT#10	XI2/XI0/XI0/ANOT#9	7.21709e-17
C152	VDD#102	XI3/XI0/XI1/net2#3	5.00211e-18
C153	VDD#14	XI0/XI1/XI4/net24#13	1.09794e-18
C154	GND#150	XI0/XI1/D#19	1.45214e-17
C155	XI3/XI1/Q#9	GND#84	1.37107e-17
C156	VDD#109	VDD	4.74455e-17
C157	VDD#160	net7#6	4.16751e-18
C158	PHI#5	XI0/XI1/Q	1.20146e-17
C159	net14#21	VDD#156	7.44569e-18
C160	RST#5	GND#138	7.22408e-18
C161	XI0/XI0/XI0/BNOT#7	XI0/XI0/XI0/ANOT#9	4.40775e-18
C162	RST#2	GND#148	6.19589e-18
C163	VDD#138	VDD	2.30186e-17
C164	GND#95	GND#72	8.36698e-18
C165	XI0/XI1/Q#7	VDD	1.11747e-17
C166	VDD#142	XI3/XI1/D#10	1.29802e-17
C167	XI3/XI1/XI4/net24#11	XI3/XI1/XI4/net24#10	7.53548e-18
C168	XI3/XI1/XI4/PHINOT#2	PHI#20	2.96218e-17
C169	XI2/XI1/XI4/net24#13	XI2/XI1/Q#7	3.21387e-18
C170	VDD#104	XI3/XI0/XI0/BNOT#3	8.47855e-18
C171	XI2/XI1/XI4/net24#9	XI2/XI1/XI4/PHINOT#3	8.28164e-18
C172	GND#78	XI3/XI1/XI4/PHINOT#3	2.02958e-18
C173	XI2/XI1/XI4/net24#11	XI2/XI1/D#4	3.45102e-18
C174	VDD#174	XI0/net1#3	2.93418e-18
C175	XI3/XI1/Q#11	SOUT3#19	7.03151e-18
C176	SOUT1#16	SOUT1#19	1.38255e-17
C177	GND#62	XI2/XI1/Q#3	4.41398e-18
C178	XI0/XI1/Q#5	VDD	1.57977e-17
C179	net21#7	XI3/XI0/XI0/BNOT#3	5.54788e-17
C180	SOUT1#20	net14#21	2.65633e-17
C181	SOUT3#11	XI3/XI0/XI0/BNOT#14	3.25292e-18
C182	XI1/XI0/XI1/net2#15	net14#15	8.93527e-18
C183	VDD#163	VDD#36	1.0238e-17
C184	GND#148	XI0/XI1/XI4/net24#3	4.14351e-18
C185	XI3/XI1/XI4/PHINOT#4	PHI#19	8.09825e-18
C186	XI2/XI0/XI0/ANOT#4	SOUT2#1	1.96312e-18
C187	GND#32	GND#141	1.0238e-17
C188	VDD#105	XI3/XI1/Q#2	2.47832e-18
C189	SOUT2	VDD#112	1.57577e-17
C190	net21#15	XI2/XI0/XI1/net2#2	3.27874e-18
C191	RST#5	XI1/net1	2.28596e-17
C192	SOUT3#14	XI3/XI1/Q	7.83548e-18
C193	RST#10	XI3/net1	3.14306e-18
C194	XI3/XI1/D#17	PHI#24	1.97458e-18
C195	GND#139	XI1/XI1/Q#9	1.24572e-17
C196	SOUT2#5	net14#5	4.43091e-17
C197	XI2/XI1/Q#9	SOUT2#19	5.37314e-18
C198	XI0/XI1/XI4/net24#6	XI0/XI1/D	1.8988e-18
C199	VDD#50	SOUT1#20	4.21807e-18
C200	XI1/XI1/D#2	XI1/XI1/XI4/PHINOT#2	1.00039e-18
C201	XI3/XI1/XI4/net24#4	PHI#24	3.61375e-17
C202	GND#84	SOUT3#16	4.02471e-17
C203	SOUT1#24	XI1/XI0/XI0/BNOT#11	2.12646e-17
C204	GND#143	XI1/XI1/XI4/PHINOT#6	1.36671e-17
C205	XI3/XI1/XI4/net24#11	VDD	4.65294e-18
C206	PHI#5	VDD#22	5.40385e-18
C207	GND#120	SOUT3#19	3.10131e-18
C208	SOUT1#8	VDD#161	5.47184e-18
C209	VDD#138	net21#6	4.16751e-18
C210	PHI#11	XI1/XI1/Q#7	3.39064e-17
C211	GND#138	GND#40	9.30871e-18
C212	GND#121	XI3/XI1/D#17	4.75796e-18
C213	VDD#131	VDD	7.55008e-17
C214	net21#19	VDD#141	1.34565e-17
C215	XI2/XI1/XI4/net24#2	XI2/XI1/Q#12	1.3891e-17
C216	XI3/net1#9	VDD	1.98755e-17
C217	GND#125	GND#70	9.24934e-18
C218	VDD#8	CIN#1	1.73636e-18
C219	PHI#23	XI3/XI1/Q#7	3.39064e-17
C220	VDD#94	VDD#93	1.68878e-17
C221	XI0/XI1/XI4/net24#12	PHI#5	4.06087e-17
C222	VDD#112	XI2/XI1/Q#3	1.24354e-18
C223	XI3/XI1/XI4/net24#9	XI3/XI1/XI4/PHINOT#2	1.74823e-18
C224	GND#138	XI1/XI0/XI1/net2	2.76367e-18
C225	XI3/XI1/D#20	PHI#23	2.73964e-17
C226	VDD#112	XI2/XI1/Q	2.29584e-18
C227	XI3/net1#4	VDD	2.62325e-17
C228	VDD#143	VDD#83	1.02424e-17
C229	XI2/XI1/XI4/PHINOT#4	PHI#13	8.09825e-18
C230	GND#114	SOUT0#10	7.13064e-18
C231	XI2/XI0/XI1/net2#15	net14#5	7.43893e-18
C232	SOUT0#16	SOUT0#18	1.30402e-17
C233	net7#10	net7#11	7.3184e-18
C234	XI2/XI1/XI4/net24#6	XI2/XI1/D#2	9.87705e-18
C235	XI3/XI0/XI0/ANOT#6	GND#72	1.48844e-17
C236	net7#21	VDD#169	6.72863e-18
C237	VDD#46	net7#6	4.0872e-18
C238	XI1/XI1/Q#6	VDD#123	1.9494e-18
C239	XI0/XI1/D#20	PHI#5	2.73964e-17
C240	net14#19	VDD#68	1.37441e-17
C241	RST#11	GND#124	6.31281e-18
C242	GND#36	XI1/XI0/XI0/ANOT#2	4.32997e-18
C243	VDD#133	XI3/XI0/XI1/net2#2	1.25381e-18
C244	XI2/XI1/Q#9	XI2/XI1/XI4/net24#3	1.58103e-18
C245	GND#109	XI1/XI0/XI0/BNOT#7	1.31853e-17
C246	GND#2	XI0/XI0/XI0/ANOT#6	4.05316e-17
C247	RST#5	GND#147	7.91186e-18
C248	VDD#172	VDD	1.44935e-17
C249	GND#70	XI3/XI1/XI4/PHINOT#6	4.0951e-17
C250	XI2/XI1/Q#7	XI2/XI1/XI4/PHINOT#2	9.18965e-19
C251	XI2/XI1/Q#5	XI2/XI1/Q#4	9.30041e-18
C252	SOUT1#20	RST#8	2.00652e-17
C253	net21#19	XI3/XI0/XI0/ANOT#2	1.52499e-17
C254	GND#22	GND#113	8.15798e-18
C255	SOUT3#20	COUT#7	2.65633e-17
C256	XI0/XI1/Q#6	VDD	9.99629e-18
C257	net7#9	SOUT1#9	3.7545e-17
C258	XI2/XI1/XI4/net24#6	XI2/XI1/XI4/net24#5	6.84508e-18
C259	XI3/XI1/Q#7	XI3/XI1/XI4/PHINOT	1.21362e-17
C260	XI3/XI0/XI0/BNOT#11	SOUT3#22	7.23396e-18
C261	XI2/XI1/XI4/PHINOT#6	XI2/XI1/XI4/PHINOT#7	4.46757e-18
C262	GND#54	GND#132	1.0238e-17
C263	XI2/XI0/XI0/ANOT	net14#7	1.29274e-18
C264	VDD#66	XI2/XI1/D#3	1.58831e-18
C265	VDD#10	XI0/net1#3	3.96888e-18
C266	XI3/XI0/XI0/BNOT#4	net21#7	2.43471e-17
C267	XI1/XI0/XI1/net2#15	net7#5	7.43893e-18
C268	VDD#98	net21#6	4.0872e-18
C269	XI1/net1#9	VDD#158	1.3419e-18
C270	XI0/XI0/XI1/net2#16	VDD	3.04753e-18
C271	GND#148	XI0/XI1/XI4/net24#4	2.22377e-18
C272	GND#26	PHI#9	5.08165e-18
C273	SOUT3#2	VDD#141	4.81645e-18
C274	XI1/XI0/XI0/ANOT#4	SOUT1#2	5.09768e-18
C275	XI2/XI1/XI4/net24	XI2/XI1/D#4	2.39789e-18
C276	XI0/XI1/Q#12	XI0/XI1/XI4/PHINOT#2	2.90831e-18
C277	XI0/XI0/XI0/ANOT#6	CIN#3	5.33566e-18
C278	XI2/XI1/XI4/net24#6	XI2/XI1/XI4/PHINOT#3	5.17189e-18
C279	XI3/XI0/XI0/ANOT#4	SOUT3#2	5.09768e-18
C280	RST#5	GND#30	1.03647e-17
C281	XI2/XI1/XI4/net24#13	PHI#17	9.76906e-18
C282	PHI#11	VDD#48	5.40385e-18
C283	XI0/XI1/D#20	VDD	3.67809e-18
C284	SOUT0#19	XI0/XI1/Q#2	6.59904e-18
C285	VDD#169	net7#10	1.49363e-17
C286	VDD#161	XI1/net1#9	1.70357e-18
C287	GND#150	XI0/XI1/D#2	3.24657e-18
C288	SOUT2#20	XI2/XI0/XI1/net2#3	1.51276e-18
C289	XI3/net1#9	net21#8	1.55592e-17
C290	GND#122	XI3/XI1/D	2.42413e-18
C291	XI0/XI1/Q#12	XI0/XI1/XI4/net24#13	1.81832e-17
C292	XI0/XI1/D#2	XI0/XI1/XI4/PHINOT#2	1.00039e-18
C293	XI1/XI1/XI4/net24#11	XI1/XI1/D#4	3.45102e-18
C294	VDD#108	VDD	8.65204e-17
C295	XI0/XI1/D#10	RST#3	3.88703e-18
C296	XI2/XI1/XI4/net24#12	PHI#17	4.06087e-17
C297	XI3/XI0/XI1/net2#13	GND#86	1.11306e-17
C298	GND#148	XI0/XI1/D#17	4.75796e-18
C299	VDD#166	XI0/XI0/XI1/net2#2	1.25381e-18
C300	VDD#159	net7#7	3.76854e-18
C301	VDD#137	VDD	2.13492e-17
C302	GND#114	SOUT0#22	9.0763e-18
C303	XI3/XI1/D#17	XI3/XI1/Q#12	5.03747e-17
C304	GND#150	XI0/XI1/XI4/net24#6	1.96676e-17
C305	GND#16	XI0/XI1/XI4/net24#3	3.76841e-18
C306	XI1/XI1/XI4/net24#12	SOUT1#14	3.08296e-18
C307	GND#123	XI3/XI1/D#2	3.24657e-18
C308	SOUT2#8	XI2/XI0/XI0/ANOT	2.40961e-17
C309	VDD#96	XI3/XI1/D#3	6.45552e-18
C310	GND#20	SOUT0#20	5.19922e-18
C311	XI3/net1#2	SOUT3#5	3.43763e-18
C312	XI3/XI1/D#6	XI3/XI1/D#5	4.49187e-18
C313	GND#4	XI0/XI1/XI4/PHINOT#6	4.0951e-17
C314	GND#62	XI2/XI1/Q#2	5.13993e-18
C315	XI1/XI1/Q#11	PHI#11	1.16343e-17
C316	XI1/XI1/D#20	XI1/XI1/D#4	9.89326e-18
C317	XI3/XI1/Q#5	XI3/XI1/XI4/PHINOT	8.79316e-18
C318	SOUT3#20	XI3/XI0/XI1/net2	2.18236e-17
C319	GND#30	XI1/XI1/D#14	2.68363e-17
C320	XI1/XI0/XI0/ANOT	net7#7	1.29274e-18
C321	XI2/XI1/D#3	PHI#16	5.34502e-17
C322	XI0/XI0/XI0/ANOT#2	CIN#8	2.9337e-18
C323	XI3/net1#9	VDD#104	2.27772e-18
C324	SOUT1#14	VDD#122	1.16528e-17
C325	VDD#142	VDD#141	1.68962e-17
C326	XI3/net1#9	XI3/XI0/XI0/BNOT#14	1.07711e-17
C327	XI3/XI1/XI4/net24#2	XI3/XI1/Q#12	1.3891e-17
C328	XI1/XI0/XI1/net2#15	SOUT1#5	5.93898e-18
C329	SOUT0#3	XI0/XI0/XI0/BNOT#2	1.91621e-18
C330	net14#17	VDD#151	6.83507e-18
C331	GND#146	XI0/XI0/XI1/net2	1.02209e-18
C332	VDD#119	GND#135	2.2414e-17
C333	VDD#104	VDD	1.04322e-17
C334	net7#15	RST#5	4.68358e-17
C335	XI1/XI1/D#6	XI1/XI1/D#5	4.49187e-18
C336	VDD#98	XI3/net1#4	3.90041e-17
C337	GND#121	net21#4	3.80483e-18
C338	VDD#130	VDD	4.74455e-17
C339	PHI#17	XI2/XI1/XI4/net24	8.89281e-18
C340	VDD#136	VDD	4.07404e-17
C341	VDD#169	XI0/XI0/XI1/net2#2	1.54384e-18
C342	VDD#70	VDD#116	1.16687e-17
C343	VDD#138	XI3/XI0/XI1/net2#15	1.7071e-18
C344	VDD#171	VDD	2.30186e-17
C345	CIN#3	SOUT0#3	7.17245e-18
C346	XI1/XI0/XI0/BNOT#10	SOUT1#2	7.16694e-18
C347	XI0/XI0/XI0/ANOT#3	CIN#9	1.57734e-18
C348	XI2/XI0/XI0/BNOT	XI2/XI0/XI0/ANOT#3	4.63673e-17
C349	net14#12	GND#138	1.3363e-17
C350	XI1/XI0/XI0/ANOT#4	VDD#165	1.1119e-17
C351	CIN#13	SOUT0#8	2.94542e-17
C352	VDD#44	XI1/XI1/D#3	6.45552e-18
C353	RST#11	XI3/net1	2.28596e-17
C354	GND#78	GND#82	1.79944e-17
C355	SOUT2#8	VDD#151	7.25049e-18
C356	SOUT1#19	SOUT1#18	3.98821e-17
C357	XI2/XI1/Q#5	VDD#117	1.53345e-17
C358	XI3/XI1/XI4/net24#9	XI3/XI1/XI4/net24#13	6.59037e-18
C359	CIN#11	XI0/net1#2	4.32779e-17
C360	RST#5	SOUT1#4	2.05565e-17
C361	XI1/XI0/XI0/ANOT#4	SOUT1#1	1.96312e-18
C362	XI0/XI1/Q#7	XI0/XI1/XI4/net24	6.2497e-18
C363	GND#6	XI0/XI0/XI0/ANOT#9	5.65589e-18
C364	XI0/XI1/D#15	XI0/XI1/D#14	4.56509e-18
C365	SOUT3#14	VDD	8.86864e-18
C366	XI3/XI1/D#10	net21#17	1.25206e-17
C367	XI3/XI0/XI1/net2#16	XI3/XI0/XI1/net2#15	7.06182e-18
C368	VDD#109	XI3/XI1/D#3	4.10481e-18
C369	XI3/XI1/XI4/net24#12	SOUT3#19	5.54297e-18
C370	XI1/XI1/XI4/PHINOT#2	XI1/XI1/XI4/net24#2	5.77081e-17
C371	COUT#1	VDD	8.95824e-18
C372	GND#137	XI1/XI0/XI1/net2	1.02209e-18
C373	XI2/XI1/XI4/net24#9	XI2/XI1/XI4/net24#2	7.14446e-18
C374	VDD#40	XI1/XI1/XI4/net24#13	1.09794e-18
C375	XI1/XI1/D#4	PHI#11	2.70764e-17
C376	XI2/XI1/D#20	XI2/XI1/XI4/net24#11	1.30924e-17
C377	PHI#4	XI0/XI1/Q	2.93097e-18
C378	GND#101	XI2/net1#16	1.74589e-17
C379	XI3/XI1/Q#5	VDD#92	6.36626e-17
C380	XI3/XI1/D#19	GND#122	1.63017e-18
C381	GND#115	GND#14	9.66245e-18
C382	XI2/XI1/D#20	XI2/XI1/D#4	9.89326e-18
C383	XI1/XI1/XI4/PHINOT#2	XI1/XI1/XI4/net24	3.28269e-17
C384	GND#74	XI3/net1	4.05515e-18
C385	XI3/XI1/Q#7	VDD#110	1.95651e-18
C386	XI3/XI0/XI0/ANOT#2	net21#8	2.9337e-18
C387	CIN#6	XI0/XI0/XI1/net2#3	1.19235e-18
C388	XI1/XI1/XI4/PHINOT#4	PHI#7	8.09825e-18
C389	XI2/XI0/XI1/net2#15	net21#15	8.93527e-18
C390	GND#52	GND#133	1.02095e-17
C391	VDD#70	XI2/XI1/XI4/net24	1.58831e-18
C392	XI0/XI1/XI4/net24#11	VDD	4.65294e-18
C393	net14#17	VDD#152	2.19992e-17
C394	SOUT3#22	VDD	9.33159e-18
C395	XI1/net1#9	XI1/XI0/XI0/BNOT#9	3.86468e-18
C396	net21#12	SOUT2#16	2.93637e-18
C397	XI2/XI1/XI4/net24#11	XI2/XI1/Q	4.03173e-18
C398	GND#78	XI3/XI1/D	3.7665e-18
C399	XI0/XI0/XI1/net2#16	SOUT0#5	2.87586e-18
C400	XI0/XI1/XI4/net24#11	PHI#5	1.50188e-17
C401	SOUT3#20	VDD	7.57963e-18
C402	XI1/XI1/D#3	PHI#10	5.34502e-17
C403	XI0/XI1/XI4/net24#13	XI0/XI1/XI4/PHINOT#2	2.64065e-17
C404	GND#22	SOUT0#10	1.12163e-17
C405	XI0/net1#9	VDD	1.98755e-17
C406	XI1/XI1/Q#9	XI1/XI1/Q#3	2.18451e-18
C407	net21#2	VDD#80	3.99391e-18
C408	XI0/net1#4	VDD	2.62325e-17
C409	XI0/XI0/XI0/BNOT#4	CIN#7	2.43471e-17
C410	COUT#7	VDD	1.1147e-17
C411	XI2/XI0/XI1/net2#16	XI2/net1#4	3.40431e-17
C412	XI2/XI0/XI0/BNOT#9	XI2/XI0/XI0/ANOT#2	4.19591e-17
C413	XI0/XI0/XI0/ANOT#9	CIN#3	1.29853e-18
C414	SOUT1#14	SOUT1#15	6.95608e-18
C415	GND#18	SOUT0#16	4.02471e-17
C416	GND#114	SOUT0#9	2.67289e-18
C417	COUT#5	VDD	1.10481e-17
C418	XI1/XI0/XI0/BNOT#9	XI1/XI0/XI0/ANOT#2	4.19591e-17
C419	VDD#136	XI3/XI0/XI1/net2#3	3.05777e-18
C420	XI0/XI1/XI4/net24#11	PHI#4	7.57347e-18
C421	XI2/XI0/XI0/ANOT#6	GND#50	1.48844e-17
C422	XI1/XI1/Q#9	GND#40	1.37107e-17
C423	GND#147	SOUT0#19	3.10131e-18
C424	XI3/XI1/D#19	PHI#21	2.62196e-18
C425	GND#92	VDD	2.72432e-17
C426	XI1/net1#9	XI1/XI0/XI0/ANOT	1.29015e-18
C427	GND#82	XI3/XI1/D#17	1.61841e-17
C428	VDD#123	XI1/XI1/D#3	4.10481e-18
C429	CIN#11	VDD#173	6.83507e-18
C430	GND#140	XI1/XI1/D#2	5.80251e-18
C431	XI1/XI1/D#16	RST#5	5.13284e-17
C432	SOUT2#24	XI2/XI0/XI0/BNOT#11	2.12646e-17
C433	XI1/XI1/D#15	net7#17	5.95074e-18
C434	GND#50	XI2/XI0/XI0/BNOT#7	4.05316e-17
C435	VDD#133	VDD	9.24489e-17
C436	PHI#17	XI2/XI1/Q#7	3.39064e-17
C437	net14#19	VDD#60	6.27963e-18
C438	XI1/net1#4	XI1/XI0/XI1/net2#3	1.41355e-18
C439	net7#21	GND#146	1.4419e-17
C440	RST#8	GND#54	1.18488e-17
C441	VDD#172	XI0/net1#9	1.70357e-18
C442	XI0/XI1/D#14	XI0/net1	2.44048e-18
C443	VDD#105	VDD	1.07942e-16
C444	GND#20	GND#147	8.84679e-18
C445	SOUT3#20	COUT#5	1.77949e-16
C446	SOUT2#10	net14#8	3.40191e-18
C447	SOUT3#22	GND#92	2.23064e-17
C448	GND#119	RST#13	2.41904e-17
C449	GND#16	XI0/XI1/XI4/net24#4	3.29561e-18
C450	VDD#104	SOUT3#22	3.78854e-17
C451	XI2/XI1/XI4/net24#11	PHI#17	1.50188e-17
C452	GND#74	GND#124	1.02095e-17
C453	GND#119	COUT#3	1.33266e-18
C454	CIN#2	VDD	2.30792e-18
C455	XI0/XI1/Q#5	XI0/XI1/XI4/net24	3.34152e-18
C456	XI3/XI0/XI0/BNOT#9	SOUT3#22	1.14498e-17
C457	XI3/XI1/XI4/net24#9	XI3/XI1/D#2	3.0624e-17
C458	XI0/XI0/XI1/net2#13	RST#2	2.21589e-17
C459	VDD#18	XI0/XI1/XI4/net24#11	6.32412e-17
C460	net21#17	VDD#141	2.19992e-17
C461	XI3/net1#9	XI3/XI0/XI0/ANOT	1.29015e-18
C462	RST#5	GND#142	6.31281e-18
C463	GND#150	GND#149	9.26445e-18
C464	XI0/XI1/Q#6	XI0/XI1/XI4/PHINOT#2	2.75539e-18
C465	VDD#166	XI0/XI0/XI1/net2	8.82071e-19
C466	XI2/XI0/XI0/ANOT#4	XI2/XI0/XI0/BNOT#10	2.24348e-18
C467	XI2/XI1/Q#11	SOUT2#19	7.03151e-18
C468	VDD#14	XI0/XI1/XI4/PHINOT	3.64808e-18
C469	PHI#2	VDD	6.36791e-17
C470	XI2/XI1/D	XI2/XI1/XI4/net24#3	2.52567e-18
C471	SOUT0#2	VDD#173	3.04495e-18
C472	SOUT0#2	VDD	9.00561e-18
C473	XI1/XI0/XI0/ANOT#4	XI1/XI0/XI0/BNOT#5	1.1098e-17
C474	GND#72	XI3/XI0/XI0/ANOT#9	5.65589e-18
C475	RST#13	COUT#3	7.49192e-18
C476	GND#32	SOUT1#4	4.09574e-18
C477	XI0/XI0/XI0/BNOT#11	SOUT0#22	7.23396e-18
C478	XI0/XI0/XI0/BNOT#7	XI0/XI0/XI0/BNOT#8	4.0203e-18
C479	XI0/XI1/XI4/net24#9	XI0/XI1/D#2	3.0624e-17
C480	VDD#112	PHI#20	2.63987e-17
C481	GND#132	GND#131	9.26445e-18
C482	XI0/net1#2	VDD	4.21525e-17
C483	XI0/XI1/XI4/PHINOT#2	XI0/XI1/XI4/net24#2	5.77081e-17
C484	XI0/XI0/XI1/net2#16	XI0/XI0/XI1/net2#15	7.06182e-18
C485	net14#2	SOUT2#2	1.06752e-17
C486	VDD#20	XI0/net1#4	3.90041e-17
C487	XI0/XI1/XI4/net24#3	PHI#6	4.68747e-17
C488	GND#120	GND#84	9.30871e-18
C489	XI1/XI1/XI4/net24#12	PHI#11	4.06087e-17
C490	XI1/XI1/D#19	XI1/XI1/XI4/PHINOT#3	2.23795e-18
C491	VDD#129	VDD	8.65204e-17
C492	VDD#171	XI0/XI0/XI1/net2#15	1.7071e-18
C493	GND#124	XI3/net1	4.15538e-18
C494	GND#121	XI3/XI1/XI4/net24#4	2.22377e-18
C495	XI1/XI1/XI4/net24#4	PHI#12	3.61375e-17
C496	XI1/XI1/Q#6	XI1/XI1/XI4/net24	1.04447e-18
C497	VDD#155	XI1/XI0/XI1/net2	8.82071e-19
C498	XI3/XI1/Q#7	XI3/XI1/XI4/net24	6.2497e-18
C499	VDD#170	VDD	2.13492e-17
C500	XI0/XI0/XI1/net2#13	GND#20	1.11306e-17
C501	PHI#6	XI0/XI1/Q#2	2.86362e-18
C502	SOUT2#8	VDD#68	1.33308e-17
C503	RST#8	XI2/net1	2.28596e-17
C504	VDD#100	SOUT3	4.09262e-18
C505	XI0/XI1/XI4/PHINOT#2	VDD	3.27746e-18
C506	SOUT3#8	VDD#94	1.33308e-17
C507	VDD#48	XI1/XI1/Q	4.68876e-18
C508	XI3/XI0/XI0/ANOT#6	SOUT3#3	2.75761e-18
C509	GND#116	SOUT0#3	5.38904e-18
C510	XI0/net1#9	XI0/XI0/XI0/BNOT#14	1.07711e-17
C511	XI1/XI1/D#17	XI1/XI1/XI4/net24#2	6.90619e-18
C512	SOUT3	VDD#108	3.91522e-17
C513	XI1/XI1/Q#6	VDD#40	1.63056e-17
C514	RST#11	SOUT3#4	2.05565e-17
C515	XI1/XI1/Q#9	XI1/XI1/Q#11	1.53602e-18
C516	XI1/XI0/XI1/net2#13	SOUT1#5	2.17512e-17
C517	SOUT1#20	net14#14	1.77949e-16
C518	VDD#141	XI3/net1#2	8.21861e-18
C519	XI1/XI0/XI1/net2#13	net14#15	8.86742e-18
C520	SOUT1#22	GND#106	2.23064e-17
C521	XI3/XI1/XI4/net24#13	XI3/XI1/XI4/PHINOT#2	2.64065e-17
C522	VDD#158	net14#10	1.49363e-17
C523	RST#5	net7#12	7.49192e-18
C524	GND#121	XI3/XI1/Q#9	1.24572e-17
C525	GND#101	GND#58	9.66245e-18
C526	SOUT0#16	XI0/XI1/Q#3	4.25775e-18
C527	XI0/net1#9	VDD#26	2.27772e-18
C528	SOUT1#10	XI1/XI0/XI0/BNOT#11	3.84272e-17
C529	XI3/XI1/D#16	XI3/XI1/D#15	9.36359e-18
C530	XI2/XI1/Q#9	PHI#18	4.56241e-18
C531	SOUT2#22	net21#21	1.19989e-16
C532	XI2/XI1/D#10	XI2/net1#2	7.8648e-18
C533	RST#5	GND#144	1.64699e-17
C534	PHI#16	XI2/XI1/Q	2.93097e-18
C535	VDD#26	VDD	1.04322e-17
C536	GND#107	SOUT1#22	9.0763e-18
C537	XI1/XI1/D#19	XI1/XI1/XI4/PHINOT#2	8.83178e-18
C538	XI0/XI0/XI0/BNOT#10	CIN#13	1.41727e-16
C539	XI1/XI0/XI0/BNOT#5	SOUT1#2	1.8238e-17
C540	GND#128	XI2/XI0/XI1/net2	1.02209e-18
C541	SOUT1#6	net7#5	3.39838e-18
C542	XI3/XI1/Q#12	XI3/XI1/D#20	2.28141e-17
C543	net14#6	XI2/XI0/XI1/net2#3	1.19235e-18
C544	SOUT2#18	XI2/XI1/Q#2	5.04785e-18
C545	VDD#169	VDD	4.07404e-17
C546	GND#42	SOUT1#20	5.19922e-18
C547	net21#17	RST#11	7.73029e-18
C548	XI3/net1#9	VDD#136	1.3419e-18
C549	XI2/XI0/XI0/BNOT#14	XI2/XI0/XI0/BNOT#4	7.00366e-18
C550	SOUT0#22	net7#21	1.19989e-16
C551	XI1/XI1/D#2	XI1/XI1/XI4/net24#2	4.04498e-17
C552	XI1/XI0/XI1/net2#13	GND#139	1.3169e-17
C553	XI3/XI1/D#14	GND#76	1.28303e-17
C554	GND#100	net14#9	4.17672e-18
C555	GND#22	SOUT0#9	5.27208e-18
C556	GND#38	XI1/XI1/Q#9	3.30192e-17
C557	XI0/XI1/D#4	VDD	8.75864e-18
C558	XI3/XI1/Q#5	XI3/XI1/XI4/net24	3.34152e-18
C559	net7#5	XI1/XI0/XI1/net2#2	4.87283e-18
C560	SOUT0#14	VDD	8.86864e-18
C561	CIN#7	XI0/XI0/XI0/BNOT#3	5.54788e-17
C562	XI3/XI0/XI1/net2#13	XI3/XI0/XI1/net2	2.66668e-18
C563	PHI#5	VDD	6.78718e-17
C564	VDD#131	XI0/XI1/XI4/PHINOT	4.411e-18
C565	XI0/XI1/XI4/net24#12	SOUT0#19	5.54297e-18
C566	net7#10	VDD	8.95824e-18
C567	GND#121	XI3/XI1/XI4/net24#3	4.14351e-18
C568	net14#17	XI2/net1#2	4.32779e-17
C569	SOUT3#14	SOUT3	3.64962e-17
C570	SOUT1#24	XI1/XI0/XI0/BNOT#9	6.98011e-18
C571	GND#139	GND#38	1.0238e-17
C572	XI2/XI1/XI4/net24#4	PHI#18	3.61375e-17
C573	XI1/XI0/XI0/BNOT#10	net7#19	1.41727e-16
C574	RST#2	CIN#4	1.53357e-17
C575	VDD#122	XI1/XI1/Q	4.97335e-18
C576	XI0/XI0/XI0/BNOT#11	CIN#9	3.59305e-18
C577	XI2/XI1/D#20	VDD#70	2.68757e-17
C578	GND#139	XI1/XI1/D#17	4.75796e-18
C579	XI0/XI0/XI1/net2#2	VDD	5.47535e-18
C580	XI1/XI1/XI4/PHINOT#9	PHI#8	1.01564e-16
C581	GND#80	XI3/XI0/XI0/ANOT#2	4.32997e-18
C582	XI3/XI1/XI4/net24#12	SOUT3#14	3.08296e-18
C583	SOUT0#22	VDD	9.33159e-18
C584	SOUT3#8	VDD#140	7.25049e-18
C585	VDD#109	PHI#22	4.96959e-18
C586	XI0/XI1/D#17	XI0/XI1/Q#12	5.03747e-17
C587	XI2/XI1/XI4/net24#6	XI2/XI1/D	1.8988e-18
C588	XI0/XI1/Q#7	XI0/XI1/XI4/PHINOT#2	9.18965e-19
C589	SOUT0#20	VDD	7.57963e-18
C590	XI0/XI0/XI0/BNOT#4	VDD	1.9561e-18
C591	XI1/XI1/D#17	XI1/XI1/Q#9	7.82323e-18
C592	SOUT1#18	PHI#11	1.77809e-17
C593	XI3/XI1/Q#6	VDD#92	1.63056e-17
C594	PHI#24	XI3/XI1/Q#2	2.86362e-18
C595	VDD#72	XI2/XI0/XI1/net2#16	1.4293e-18
C596	VDD#137	VDD#136	1.8229e-17
C597	SOUT1#22	net7#8	5.05993e-18
C598	GND#26	XI1/XI1/XI4/PHINOT#6	4.0951e-17
C599	GND#141	SOUT1#4	3.19662e-18
C600	XI3/XI1/XI4/net24#6	XI3/XI1/D#2	9.87705e-18
C601	XI3/XI0/XI0/ANOT#9	SOUT3#3	2.35212e-17
C602	net7#21	VDD	1.1147e-17
C603	GND#92	VDD#134	1.53265e-17
C604	net14#8	XI2/XI0/XI0/BNOT#4	3.19507e-18
C605	XI0/XI1/D#19	XI0/XI1/XI4/net24#9	4.55106e-18
C606	XI3/XI1/D#15	net21#17	5.95074e-18
C607	GND#34	XI1/XI1/D#2	9.24969e-18
C608	GND#93	SOUT3#10	7.13064e-18
C609	net7#14	VDD	1.10481e-17
C610	RST#8	GND#132	9.12929e-18
C611	GND#148	PHI#6	5.83194e-18
C612	PHI#8	VDD	1.10308e-16
C613	XI0/XI1/XI4/PHINOT#2	XI0/XI1/XI4/net24	3.28269e-17
C614	VDD#105	XI3/XI1/Q#3	1.24354e-18
C615	XI3/XI1/Q#5	VDD#110	1.53345e-17
C616	RST#5	XI1/XI1/D#6	1.04408e-17
C617	GND#113	VDD	2.72001e-17
C618	SOUT1#2	VDD	9.00561e-18
C619	VDD#42	SOUT1#7	8.24977e-18
C620	GND#129	XI2/XI0/XI1/net2	2.76367e-18
C621	XI0/XI1/D#2	XI0/XI1/XI4/PHINOT#3	3.94365e-17
C622	VDD#92	XI3/XI1/XI4/PHINOT	3.64808e-18
C623	XI3/XI1/D#19	GND#78	2.48425e-18
C624	GND#128	VDD#144	7.65081e-17
C625	XI1/net1#2	VDD	4.21525e-17
C626	GND#28	XI1/XI0/XI0/BNOT#7	4.05316e-17
C627	RST#1	XI0/net1	3.14306e-18
C628	XI0/XI0/XI0/BNOT#10	XI0/XI0/XI0/ANOT#9	7.21709e-17
C629	XI3/XI1/XI4/PHINOT#9	PHI#20	1.01564e-16
C630	VDD#166	VDD	7.78897e-17
C631	SOUT0#10	XI0/XI0/XI0/BNOT#11	3.84272e-17
C632	VDD#52	XI1/XI0/XI0/BNOT#4	1.39714e-18
C633	XI2/XI1/Q#11	PHI#18	1.32498e-17
C634	GND#82	XI3/XI1/XI4/net24#4	3.29561e-18
C635	XI1/XI0/XI0/BNOT#7	SOUT1#3	5.63912e-18
C636	PHI#10	XI1/XI1/Q	2.93097e-18
C637	SOUT0#19	SOUT0#18	3.98821e-17
C638	GND#58	XI2/XI0/XI0/ANOT#2	4.32997e-18
C639	GND#6	SOUT0#3	4.36955e-18
C640	VDD#144	XI2/XI0/XI1/net2	8.82071e-19
C641	VDD#126	VDD	9.39951e-17
C642	GND#12	GND#16	1.79944e-17
C643	COUT#1	XI3/XI0/XI1/net2#3	6.65581e-18
C644	SOUT3	VDD#105	1.57577e-17
C645	net7#6	XI1/XI0/XI1/net2#3	1.19235e-18
C646	XI1/XI1/XI4/PHINOT#2	VDD	3.27746e-18
C647	PHI#14	VDD#56	6.00445e-18
C648	XI2/XI0/XI0/ANOT#9	net14#2	4.97779e-17
C649	SOUT3#8	VDD#139	5.47184e-18
C650	VDD#72	XI2/XI0/XI1/net2#3	1.01229e-18
C651	XI2/XI0/XI0/BNOT#14	net14#7	1.32694e-17
C652	XI1/XI0/XI0/ANOT#4	VDD#34	2.2775e-17
C653	COUT#3	SOUT3#16	2.93637e-18
C654	XI2/XI0/XI1/net2#2	SOUT2#20	1.29961e-17
C655	net14#17	VDD#64	1.45914e-17
C656	SOUT0#19	XI0/XI1/Q#3	5.30351e-18
C657	XI1/XI1/XI4/net24#11	SOUT1#14	9.24112e-18
C658	GND#137	VDD#155	7.65081e-17
C659	XI3/XI0/XI0/BNOT#14	SOUT3#22	8.52113e-18
C660	SOUT2#8	VDD#150	5.47184e-18
C661	SOUT3#14	PHI#23	1.23563e-17
C662	XI1/XI1/XI4/net24#11	PHI#11	1.50188e-17
C663	XI2/XI0/XI1/net2#13	net21#15	8.86742e-18
C664	VDD#28	VDD	1.49508e-17
C665	RST#8	SOUT2#4	2.05565e-17
C666	GND#131	GND#56	1.01892e-17
C667	net14#7	XI2/XI0/XI0/BNOT#3	5.54788e-17
C668	VDD#162	SOUT1#6	4.21273e-18
C669	GND#108	XI1/XI0/XI0/BNOT	2.7139e-18
C670	XI3/XI1/Q#7	XI3/XI1/XI4/PHINOT#2	9.18965e-19
C671	GND#82	XI3/XI1/XI4/net24#3	3.76841e-18
C672	VDD#88	XI3/net1#2	1.39754e-17
C673	XI1/XI1/XI4/net24#13	XI1/XI1/Q#7	3.21387e-18
C674	CIN#2	VDD#1	2.42465e-18
C675	XI0/XI0/XI0/ANOT#4	SOUT0#1	1.96312e-18
C676	XI2/XI0/XI0/BNOT#2	XI2/XI0/XI0/ANOT#2	6.90696e-17
C677	VDD#165	VDD	7.27918e-17
C678	XI0/XI1/XI4/net24#6	XI0/XI1/D#2	9.87705e-18
C679	XI3/XI1/D#4	PHI#23	2.70764e-17
C680	XI0/XI1/D#2	XI0/XI1/XI4/net24#2	4.04498e-17
C681	XI0/XI1/XI4/PHINOT#4	PHI#1	8.09825e-18
C682	XI2/XI1/D#2	XI2/XI1/XI4/net24#4	1.54296e-18
C683	XI2/XI0/XI1/net2#13	GND#64	1.11306e-17
C684	GND#4	PHI#3	5.08165e-18
C685	SOUT2#20	VDD#147	2.36869e-17
C686	XI0/XI0/XI0/ANOT#9	SOUT0#2	2.69483e-18
C687	GND#139	net7#4	3.80483e-18
C688	XI2/XI1/Q#9	XI2/XI1/Q#11	1.53602e-18
C689	XI2/XI1/D#20	PHI#17	2.73964e-17
C690	XI1/XI1/D#17	PHI#12	1.97458e-18
C691	VDD#110	XI3/XI1/XI4/PHINOT	4.411e-18
C692	XI2/XI0/XI0/BNOT#11	XI2/XI0/XI0/BNOT#9	1.98917e-17
C693	XI1/XI1/D#20	PHI#11	2.73964e-17
C694	XI1/net1#9	VDD#159	7.01142e-18
C695	GND#12	XI0/XI1/XI4/PHINOT#3	2.02958e-18
C696	XI1/net1	SOUT1#5	4.53739e-18
C697	XI2/XI1/D#15	XI2/net1#2	3.59645e-18
C698	XI0/XI1/D#4	PHI#5	2.70764e-17
C699	XI3/XI1/D#14	RST#11	5.02859e-17
C700	VDD#52	net7#7	4.04071e-18
C701	XI3/XI1/XI4/net24#9	XI3/XI1/XI4/net24#2	7.14446e-18
C702	net14#10	SOUT1#20	4.66076e-17
C703	XI2/XI1/XI4/net24#9	XI2/XI1/Q#12	4.7443e-18
C704	XI2/XI1/XI4/net24#13	XI2/XI1/XI4/net24#2	1.71266e-17
C705	XI1/XI1/D#4	VDD	8.75864e-18
C706	GND#152	GND#4	9.24934e-18
C707	SOUT0#11	XI0/XI0/XI0/ANOT	8.09714e-18
C708	SOUT1#14	SOUT1#18	1.77557e-17
C709	XI2/net1#9	VDD#78	2.27772e-18
C710	VDD#88	net21#17	2.54235e-17
C711	GND#107	SOUT1#9	2.67289e-18
C712	VDD#30	VDD	1.68456e-17
C713	VDD#161	SOUT1#7	2.63522e-18
C714	PHI#11	VDD	6.78718e-17
C715	VDD#56	XI2/XI1/XI4/PHINOT#4	5.55471e-17
C716	VDD#176	VDD#5	1.02424e-17
C717	VDD#62	net14#17	2.54235e-17
C718	SOUT1#2	VDD#163	4.81645e-18
C719	VDD#125	VDD	1.32558e-16
C720	XI3/XI0/XI0/BNOT#9	net21#19	1.54043e-17
C721	XI1/XI1/D#14	GND#142	6.94823e-18
C722	XI2/XI1/XI4/net24#11	VDD#74	1.81691e-17
C723	GND#20	XI0/XI0/XI1/net2	4.49691e-18
C724	XI2/XI0/XI1/net2#16	XI2/XI0/XI1/net2#15	7.06182e-18
C725	XI2/XI0/XI1/net2#13	GND#130	1.3169e-17
C726	VDD#31	VDD	2.12045e-17
C727	GND#8	XI0/XI1/D#14	2.68363e-17
C728	SOUT0#24	XI0/XI0/XI0/BNOT#2	5.12165e-17
C729	XI2/XI1/D#2	XI2/XI1/D#17	3.60142e-18
C730	XI1/XI1/D#15	RST#5	4.36037e-17
C731	XI2/XI1/Q#11	XI2/XI1/Q#2	3.35663e-18
C732	XI2/XI0/XI0/BNOT#10	net14#2	2.58085e-18
C733	XI1/XI0/XI1/net2#2	VDD	5.47535e-18
C734	GND#120	XI3/XI1/Q#3	2.16945e-18
C735	XI3/net1#2	SOUT3#6	1.96305e-17
C736	XI3/net1#4	net21#6	1.35025e-17
C737	SOUT0#18	PHI#5	1.77809e-17
C738	GND#54	GND#53	7.9864e-18
C739	net7#19	VDD#42	1.37441e-17
C740	GND#82	XI3/XI1/Q#9	3.30192e-17
C741	SOUT2#24	XI2/XI0/XI0/BNOT#9	6.98011e-18
C742	XI1/XI0/XI0/ANOT#4	VDD	9.31981e-18
C743	net14#14	RST#8	4.02246e-17
C744	XI1/XI0/XI0/BNOT#4	VDD	1.9561e-18
C745	XI2/XI1/XI4/net24#12	SOUT2#19	5.54297e-18
C746	VDD#86	SOUT3#1	4.22292e-18
C747	SOUT2#2	VDD#151	3.04495e-18
C748	GND#16	XI0/XI1/D#17	1.61841e-17
C749	VDD#38	SOUT1#6	4.07255e-18
C750	GND#50	XI2/XI0/XI0/ANOT#9	5.65589e-18
C751	VDD#80	XI3/XI0/XI0/ANOT#4	5.51165e-17
C752	XI1/net1#9	XI1/XI0/XI0/BNOT#14	1.07711e-17
C753	GND#88	SOUT3#10	1.12163e-17
C754	VDD#153	net14#19	3.06108e-18
C755	GND#94	XI3/net1#16	1.74589e-17
C756	XI3/XI1/Q#6	XI3/XI1/D#20	8.17481e-17
C757	VDD#2	CIN#1	5.53658e-18
C758	XI0/XI1/XI4/net24#2	XI0/XI1/XI4/PHINOT#3	1.97764e-17
C759	PHI#14	VDD	1.10308e-16
C760	PHI#8	XI1/XI1/XI4/PHINOT#4	4.3751e-18
C761	SOUT2#10	SOUT2#22	5.91301e-18
C762	XI1/XI1/XI4/PHINOT#9	VDD	4.78049e-18
C763	SOUT2#11	XI2/XI0/XI0/ANOT	8.09714e-18
C764	SOUT2#2	VDD	9.00561e-18
C765	XI0/XI1/D#16	RST#2	5.30268e-17
C766	XI1/XI1/XI4/PHINOT#4	VDD	2.14306e-17
C767	VDD#26	VDD#169	1.09613e-17
C768	XI3/XI1/XI4/net24#11	XI3/XI1/D#3	3.27281e-18
C769	VDD#78	VDD#77	1.35961e-17
C770	XI3/XI1/XI4/PHINOT#6	PHI#21	9.47309e-18
C771	XI2/net1#2	VDD	4.21525e-17
C772	XI3/net1	SOUT3#5	4.53739e-18
C773	XI1/XI1/D#10	VDD	1.26139e-17
C774	VDD#78	VDD#147	1.09613e-17
C775	net14#10	XI1/XI0/XI1/net2#2	5.88268e-18
C776	XI2/XI1/Q#7	XI2/XI1/Q#5	9.68451e-18
C777	XI2/XI0/XI0/ANOT#6	SOUT2#3	2.75761e-18
C778	SOUT0#22	CIN#8	5.05993e-18
C779	PHI#20	XI3/XI1/XI4/PHINOT#4	4.3751e-18
C780	VDD#24	net7#10	5.51165e-17
C781	XI3/XI1/XI4/net24#11	SOUT3#14	9.24112e-18
C782	VDD#140	VDD#90	1.0238e-17
C783	GND#121	PHI#24	5.83194e-18
C784	XI2/XI1/XI4/PHINOT#2	VDD	3.27746e-18
C785	GND#36	XI1/XI0/XI0/BNOT	4.9463e-18
C786	VDD#28	net7	5.53658e-18
C787	SOUT1#20	RST#5	1.76518e-17
C788	VDD#76	net21#10	5.51165e-17
C789	net7#7	XI1/XI0/XI0/BNOT#3	5.54788e-17
C790	SOUT2#20	net21#21	2.65633e-17
C791	XI3/net1#16	SOUT3#10	4.33498e-18
C792	GND#93	GND#88	9.65661e-18
C793	XI2/XI0/XI0/ANOT#4	XI2/XI0/XI0/BNOT#5	1.1098e-17
C794	GND#148	GND#16	1.0238e-17
C795	RST#5	GND#143	1.95518e-17
C796	VDD#123	PHI#10	4.96959e-18
C797	SOUT0#6	CIN#5	3.39838e-18
C798	XI1/XI0/XI0/BNOT#4	VDD#158	2.37247e-18
C799	XI2/XI0/XI1/net2#15	SOUT2#5	5.93898e-18
C800	GND#139	XI1/XI1/XI4/net24#4	2.22377e-18
C801	GND#52	GND#51	7.83801e-18
C802	XI3/XI1/D#14	XI3/net1	2.44048e-18
C803	CIN#13	VDD#8	6.30034e-18
C804	GND#119	XI3/XI0/XI1/net2	1.0422e-18
C805	net14#2	XI2/XI0/XI0/ANOT#4	3.09365e-18
C806	VDD#92	VDD#96	3.93119e-17
C807	XI3/XI0/XI1/net2#15	SOUT3#5	5.93898e-18
C808	VDD#164	VDD	1.8633e-17
C809	RST#8	XI2/net1#2	3.74826e-18
C810	net21#12	net21#13	4.31453e-18
C811	VDD#100	SOUT3#14	5.47763e-17
C812	CIN#13	XI0/XI0/XI0/ANOT#2	1.52499e-17
C813	XI0/XI1/D#16	XI0/XI1/D#15	9.36359e-18
C814	RST#8	GND#129	7.22408e-18
C815	net21#5	XI3/XI0/XI1/net2#2	4.87283e-18
C816	XI0/XI1/XI4/net24#4	XI0/XI1/Q#12	2.8824e-17
C817	VDD#40	VDD#124	1.16687e-17
C818	net7#17	RST#5	7.73029e-18
C819	GND#44	SOUT1#9	5.27208e-18
C820	CIN#11	SOUT0#5	2.7909e-17
C821	GND#40	XI1/XI1/Q#2	5.13993e-18
C822	XI0/XI1/D#17	XI0/XI1/Q#9	7.82323e-18
C823	SOUT0#14	XI0/XI1/Q	7.83548e-18
C824	XI3/XI1/Q#6	VDD#110	4.14214e-18
C825	GND#84	XI3/XI1/Q#3	4.41398e-18
C826	GND#147	SOUT0#18	1.34133e-17
C827	XI2/XI1/XI4/net24#2	XI2/XI1/XI4/net24#4	1.52005e-18
C828	VDD#104	VDD#103	1.35961e-17
C829	VDD#136	XI3/XI0/XI1/net2#2	1.54384e-18
C830	XI0/XI1/D#15	XI0/net1	1.96101e-17
C831	SOUT1#16	XI1/XI1/Q#3	4.25775e-18
C832	GND#109	GND#28	8.36698e-18
C833	XI3/XI1/D#15	RST#11	4.36037e-17
C834	RST#8	GND#42	1.13456e-17
C835	GND#129	SOUT2#18	1.34133e-17
C836	VDD#164	XI1/XI1/D#10	1.29802e-17
C837	XI1/XI1/D#15	XI1/XI1/D#14	4.56509e-18
C838	CIN#1	SOUT0#1	3.65393e-18
C839	PHI#17	XI2/XI1/XI4/PHINOT#2	4.78246e-17
C840	XI1/XI1/D#14	GND#32	1.28303e-17
C841	XI2/XI0/XI0/BNOT#5	XI2/XI0/XI0/BNOT#6	8.47836e-18
C842	XI2/XI0/XI1/net2#13	net14#4	2.31785e-18
C843	net21#21	VDD#145	7.44569e-18
C844	XI2/XI1/D#4	VDD	8.75864e-18
C845	SOUT3#20	GND#119	1.26093e-17
C846	GND#122	GND#78	1.01892e-17
C847	XI1/XI1/Q#7	XI1/XI1/Q#6	6.45394e-18
C848	XI3/XI1/D#2	XI3/XI1/D#17	3.60142e-18
C849	XI1/XI0/XI0/BNOT#5	VDD	8.81368e-18
C850	PHI#17	VDD	6.78718e-17
C851	GND#148	XI0/XI1/Q#9	1.24572e-17
C852	SOUT3#20	VDD#136	2.36869e-17
C853	VDD#163	VDD	1.94359e-17
C854	SOUT0#16	SOUT0#17	4.09771e-18
C855	VDD#176	CIN#1	2.66145e-18
C856	VDD#105	XI3/XI1/Q	2.29584e-18
C857	VDD#92	XI3/XI1/XI4/net24	6.41722e-18
C858	net7#14	GND#146	1.08364e-16
C859	SOUT3#20	XI3/XI0/XI1/net2#3	1.51276e-18
C860	XI3/XI1/D#15	XI3/XI1/D#14	4.56509e-18
C861	SOUT0#18	VDD#126	2.18537e-17
C862	XI0/XI0/XI1/net2#16	SOUT0#6	5.16806e-18
C863	XI3/net1#4	XI3/XI0/XI1/net2#2	9.28475e-19
C864	XI3/XI0/XI0/BNOT#11	net21#8	1.64202e-18
C865	VDD#167	VDD	4.3336e-17
C866	XI0/XI0/XI0/ANOT#4	SOUT0#2	5.09768e-18
C867	GND#115	XI0/XI0/XI0/BNOT#2	3.63595e-18
C868	GND#18	XI0/XI1/Q#2	5.13993e-18
C869	XI1/net1#4	net7#6	1.35025e-17
C870	XI2/XI0/XI1/net2#2	VDD	5.47535e-18
C871	XI1/XI0/XI1/net2#13	net14#12	3.2914e-18
C872	VDD#127	VDD	5.73405e-17
C873	net21#19	SOUT3#2	6.17276e-17
C874	SOUT0#20	RST#5	2.00652e-17
C875	COUT#1	COUT#2	7.3184e-18
C876	XI2/XI1/XI4/net24#12	XI2/XI1/Q#2	2.89847e-18
C877	XI2/XI1/D#20	VDD#116	2.76988e-18
C878	XI2/XI1/D#6	GND#134	1.65584e-17
C879	GND#130	XI2/XI1/XI4/net24#4	2.22377e-18
C880	XI1/XI1/Q#6	VDD#124	4.14214e-18
C881	CIN#5	XI0/XI0/XI1/net2#2	4.87283e-18
C882	XI3/XI1/XI4/PHINOT#9	PHI#21	1.27134e-18
C883	PHI#6	XI0/XI1/Q#3	3.05252e-18
C884	net14#17	SOUT2#5	2.7909e-17
C885	XI3/XI1/XI4/net24#9	XI3/XI1/Q#12	4.7443e-18
C886	XI1/net1#9	VDD#160	3.67621e-17
C887	net7#19	VDD	7.38122e-18
C888	XI3/XI1/D#20	VDD#96	2.68757e-17
C889	XI2/XI1/Q#7	XI2/XI1/XI4/PHINOT	1.21362e-17
C890	XI2/XI0/XI0/BNOT#4	VDD	1.9561e-18
C891	RST#13	GND#86	1.13456e-17
C892	PHI#11	XI1/XI1/Q#2	2.73644e-17
C893	net7#17	VDD	6.33291e-18
C894	XI0/XI1/XI4/net24#11	VDD#130	1.56401e-17
C895	VDD#26	XI0/XI0/XI0/BNOT#3	8.47855e-18
C896	SOUT0#22	CIN#9	1.80819e-18
C897	XI1/XI1/D#6	GND#143	1.65584e-17
C898	XI0/XI0/XI0/BNOT#9	SOUT0#22	1.14498e-17
C899	GND#103	XI2/XI0/XI0/ANOT#6	1.31853e-17
C900	CIN#11	VDD#12	1.45914e-17
C901	GND#147	GND#18	9.30871e-18
C902	XI2/XI0/XI0/ANOT#9	SOUT2#3	2.35212e-17
C903	XI0/XI0/XI0/ANOT#9	CIN#13	7.0373e-18
C904	VDD#98	XI3/XI0/XI1/net2#16	1.4293e-18
C905	SOUT1#5	net7#5	4.43091e-17
C906	XI0/XI1/Q#11	XI0/XI1/Q#2	3.35663e-18
C907	PHI#20	VDD	1.10308e-16
C908	VDD#133	XI3/XI0/XI1/net2	8.86371e-19
C909	XI0/XI1/Q#7	XI0/XI1/Q#5	9.68451e-18
C910	XI3/XI1/D#2	XI3/XI1/XI4/PHINOT#2	1.00039e-18
C911	VDD#162	VDD	2.56909e-17
C912	VDD#160	VDD#46	1.0238e-17
C913	XI1/XI0/XI0/ANOT#2	XI1/XI0/XI0/BNOT#10	7.01434e-17
C914	GND#110	XI1/XI0/XI0/ANOT#6	1.31853e-17
C915	SOUT3#2	VDD	9.00561e-18
C916	SOUT3#19	XI3/XI1/Q#2	6.59904e-18
C917	XI2/XI1/D#19	PHI#15	2.62196e-18
C918	VDD#60	SOUT2#1	4.22292e-18
C919	XI1/XI1/D#19	XI1/XI1/D#2	1.57987e-18
C920	VDD#110	XI3/XI1/XI4/net24	4.3074e-18
C921	XI2/XI0/XI0/ANOT#3	net14#9	1.57734e-18
C922	VDD#14	XI0/XI1/XI4/net24	6.41722e-18
C923	XI3/net1#2	VDD	4.21525e-17
C924	net14	SOUT2#2	2.69766e-18
C925	XI2/XI1/Q#12	XI2/XI1/XI4/net24#12	1.90043e-17
C926	XI0/XI0/XI1/net2#16	CIN#5	2.63779e-17
C927	VDD#68	VDD#67	1.68878e-17
C928	GND#129	GND#62	9.30871e-18
C929	VDD#173	XI0/net1#2	9.35443e-18
C930	GND#42	XI1/XI0/XI1/net2	4.49691e-18
C931	XI3/XI1/XI4/PHINOT#2	VDD	3.27746e-18
C932	XI0/XI1/XI4/net24#9	XI0/XI1/XI4/net24#2	7.14446e-18
C933	XI0/XI0/XI1/net2#15	net7#10	6.82353e-18
C934	XI1/net1#16	SOUT1#24	5.33627e-17
C935	SOUT3#10	net21#9	4.46078e-17
C936	GND#130	XI2/XI1/Q#9	1.24572e-17
C937	GND#94	XI3/XI0/XI0/BNOT	2.7139e-18
C938	SOUT0#10	CIN#9	4.46078e-17
C939	VDD#54	net14	5.53658e-18
C940	VDD#133	GND#118	1.39542e-17
C941	XI0/net1#9	VDD#170	7.01142e-18
C942	XI2/XI0/XI1/net2#13	net21#12	3.2914e-18
C943	XI3/XI0/XI1/net2#16	SOUT3#6	5.16806e-18
C944	net14#15	XI1/XI0/XI1/net2#2	3.27874e-18
C945	VDD#138	VDD#98	1.0238e-17
C946	GND#38	XI1/XI1/D#17	1.61841e-17
C947	SOUT1#19	XI1/XI1/Q#3	5.30351e-18
C948	XI2/XI1/Q#5	XI2/XI1/XI4/PHINOT	8.79316e-18
C949	XI0/net1#9	VDD#169	1.3419e-18
C950	SOUT0#20	net7#21	2.65633e-17
C951	XI1/XI1/Q#7	VDD	1.11747e-17
C952	XI2/net1	SOUT2#5	4.53739e-18
C953	XI1/XI0/XI0/BNOT#5	net7#19	4.10074e-17
C954	XI3/XI0/XI1/net2#13	SOUT3#5	2.17512e-17
C955	RST#2	XI0/XI1/D#6	1.04408e-17
C956	XI3/XI0/XI0/BNOT#11	XI3/XI0/XI0/BNOT#9	1.98917e-17
C957	VDD#24	XI0/XI0/XI1/net2#3	5.00211e-18
C958	GND#52	XI2/net1	4.05515e-18
C959	XI1/XI1/D#17	XI1/XI1/Q#11	1.88867e-17
C960	XI1/XI1/Q#5	VDD	1.57977e-17
C961	XI2/XI0/XI1/net2#13	SOUT2#5	2.17512e-17
C962	GND#38	XI1/XI1/XI4/net24#4	3.29561e-18
C963	CIN#2	SOUT0#2	1.06752e-17
C964	XI3/net1#16	SOUT3#24	5.33627e-17
C965	XI3/XI1/D#16	RST#11	5.13284e-17
C966	PHI#12	XI1/XI1/Q#2	2.86362e-18
C967	XI2/net1#9	VDD#149	3.67621e-17
C968	SOUT2#5	RST#8	3.79452e-17
C969	RST#2	GND#8	1.03647e-17
C970	XI3/XI0/XI0/ANOT#4	VDD#86	2.2775e-17
C971	XI3/XI0/XI0/ANOT#9	net21#19	6.99675e-18
C972	XI3/XI1/XI4/net24#11	PHI#22	7.57347e-18
C973	XI2/net1#9	VDD#147	1.3419e-18
C974	XI3/XI1/D#4	VDD	8.75864e-18
C975	GND#141	XI1/XI1/XI4/PHINOT#3	3.59673e-18
C976	net21#10	net21#11	7.3184e-18
C977	XI3/XI1/XI4/net24#11	VDD#100	1.81691e-17
C978	XI3/XI1/XI4/net24#13	XI3/XI1/XI4/net24#2	1.71266e-17
C979	XI1/XI1/XI4/net24#11	XI1/XI1/D#3	3.27281e-18
C980	XI0/XI0/XI0/BNOT#5	CIN#13	4.10074e-17
C981	XI0/XI0/XI0/BNOT#9	CIN#13	1.53223e-17
C982	XI1/XI1/XI4/PHINOT#3	XI1/XI1/D	3.80638e-17
C983	PHI#23	VDD	5.43061e-17
C984	XI0/XI1/XI4/net24#12	SOUT0#14	3.08296e-18
C985	VDD#42	XI1/XI0/XI0/ANOT	4.13602e-18
C986	XI1/XI1/D#14	RST#5	5.02859e-17
C987	XI3/XI1/D#4	VDD#96	4.83878e-18
C988	VDD#26	XI0/XI0/XI0/BNOT#4	1.39714e-18
C989	XI3/XI0/XI1/net2#15	XI3/XI0/XI1/net2#2	6.41939e-18
C990	GND#149	XI0/XI1/D	2.42413e-18
C991	VDD#124	VDD	8.4118e-17
C992	XI3/XI0/XI0/BNOT#9	net21#8	9.80156e-17
C993	net7#2	SOUT1#2	1.06752e-17
C994	XI3/XI0/XI0/ANOT#4	VDD#143	1.1119e-17
C995	XI0/XI1/D#14	SOUT0#5	7.88532e-18
C996	VDD#131	XI0/XI1/XI4/net24	4.3074e-18
C997	PHI#18	XI2/XI1/Q#2	2.86362e-18
C998	XI1/XI1/Q#5	XI1/XI1/Q#4	9.30041e-18
C999	VDD#82	XI3/XI1/XI4/PHINOT#4	5.55471e-17
C1000	SOUT3#11	net21#8	1.51116e-17
C1001	SOUT3#14	VDD#108	1.16528e-17
C1002	XI3/XI0/XI1/net2#2	VDD	5.47535e-18
C1003	XI2/XI1/D#17	XI2/XI1/XI4/net24#2	6.90619e-18
C1004	GND#66	GND#65	7.74457e-18
C1005	XI3/XI1/XI4/PHINOT#3	XI3/XI1/D	3.80638e-17
C1006	SOUT1#3	XI1/XI0/XI0/BNOT#2	1.91621e-18
C1007	XI2/XI1/XI4/net24#3	PHI#18	4.68747e-17
C1008	XI1/XI1/D#16	XI1/XI1/D#15	9.36359e-18
C1009	RST#3	XI0/net1#3	2.67237e-18
C1010	GND#123	XI3/XI1/D#19	1.45214e-17
C1011	XI2/XI1/XI4/net24#12	SOUT2#14	3.08296e-18
C1012	XI3/XI0/XI0/BNOT#4	VDD	1.9561e-18
C1013	XI2/XI1/XI4/PHINOT#4	VDD#118	1.16528e-17
C1014	XI0/XI1/Q#12	XI0/XI1/D#20	2.28141e-17
C1015	VDD#161	VDD	1.44935e-17
C1016	SOUT2#22	XI2/XI0/XI0/BNOT#4	3.05405e-18
C1017	GND#60	XI2/XI1/XI4/net24#4	3.29561e-18
C1018	XI2/XI1/XI4/PHINOT#6	PHI#15	9.47309e-18
C1019	GND#92	COUT#7	9.41186e-17
C1020	SOUT3#18	GND#119	3.44305e-17
C1021	net14#15	SOUT1#20	8.75531e-17
C1022	XI1/XI1/D#17	XI1/XI1/XI4/PHINOT#3	8.962e-19
C1023	XI1/XI1/XI4/net24	XI1/XI1/D#4	2.39789e-18
C1024	XI1/net1#4	VDD#159	1.37422e-18
C1025	XI1/XI1/Q#11	XI1/XI1/Q#2	3.35663e-18
C1026	COUT#3	GND#120	1.3363e-17
C1027	GND#108	XI1/XI0/XI0/ANOT#3	4.34667e-18
C1028	GND#80	XI3/XI0/XI0/BNOT	4.9463e-18
C1029	XI2/XI1/D#14	SOUT2#5	7.88532e-18
C1030	GND#139	XI1/XI1/XI4/net24#3	4.14351e-18
C1031	XI1/XI1/XI4/PHINOT#6	XI1/XI1/XI4/PHINOT#7	4.46757e-18
C1032	XI0/XI1/Q#5	VDD#14	6.36626e-17
C1033	XI1/XI1/Q#6	VDD	9.99629e-18
C1034	VDD#8	XI0/XI0/XI0/BNOT#5	5.45774e-17
C1035	net7#10	SOUT0#20	4.66076e-17
C1036	VDD#94	VDD#139	1.0979e-17
C1037	SOUT3#3	XI3/XI0/XI0/BNOT#2	1.91621e-18
C1038	XI0/XI1/Q#7	VDD#131	1.95651e-18
C1039	SOUT0#14	SOUT0#18	1.77557e-17
C1040	XI1/XI0/XI0/BNOT#5	XI1/XI0/XI0/BNOT#6	8.47836e-18
C1041	SOUT0#5	CIN#5	4.43091e-17
C1042	GND#14	XI0/XI0/XI0/BNOT#2	1.48416e-18
C1043	XI2/net1#9	net14#8	1.55592e-17
C1044	VDD#151	XI2/net1#2	9.35443e-18
C1045	GND#141	GND#140	9.26445e-18
C1046	SOUT1#8	XI1/XI0/XI0/ANOT	2.40961e-17
C1047	XI3/XI1/XI4/PHINOT#2	XI3/XI1/XI4/net24#2	5.77081e-17
C1048	XI2/XI1/D#4	PHI#16	1.07136e-17
C1049	XI2/XI0/XI0/BNOT#5	VDD#152	1.54612e-17
C1050	VDD#148	XI2/XI0/XI1/net2#2	4.26212e-18
C1051	XI1/XI0/XI1/net2#16	VDD	3.04753e-18
C1052	SOUT2#20	net21#14	1.77949e-16
C1053	XI0/XI1/D#19	XI0/XI1/XI4/net24#6	1.52492e-17
C1054	SOUT2#10	XI2/XI0/XI0/BNOT#4	2.61929e-18
C1055	SOUT2#22	GND#99	2.23064e-17
C1056	GND#103	net14#3	3.66677e-18
C1057	GND#137	RST#8	2.41904e-17
C1058	net7#10	XI0/XI0/XI1/net2#2	5.88268e-18
C1059	XI3/XI1/XI4/net24#13	XI3/XI1/Q#7	3.21387e-18
C1060	XI3/XI1/D#17	XI3/XI1/XI4/net24#2	6.90619e-18
C1061	XI0/XI1/D#4	VDD#18	4.83878e-18
C1062	GND#122	XI3/XI1/D#17	1.58396e-18
C1063	VDD#105	PHI#25	2.49545e-17
C1064	VDD#161	XI1/XI0/XI0/ANOT	1.82797e-18
C1065	GND#133	XI2/net1	4.15538e-18
C1066	GND#102	GND#50	8.36698e-18
C1067	GND#56	XI2/XI1/XI4/PHINOT#3	2.02958e-18
C1068	XI1/XI1/D#20	VDD	3.67809e-18
C1069	XI0/XI1/XI4/net24#12	XI0/XI1/Q#2	2.89847e-18
C1070	XI0/XI1/Q#9	XI0/XI1/Q#8	3.3441e-18
C1071	VDD#153	XI2/XI1/D#10	1.29802e-17
C1072	net21#19	VDD#86	6.27963e-18
C1073	VDD#156	VDD	4.3336e-17
C1074	VDD#120	VDD	5.73405e-17
C1075	XI0/XI0/XI0/ANOT#4	XI0/XI0/XI0/BNOT#10	2.24348e-18
C1076	VDD#104	XI3/XI0/XI0/BNOT#4	1.39714e-18
C1077	CIN#11	SOUT0#6	1.79032e-18
C1078	XI1/XI1/D#19	GND#142	3.09843e-17
C1079	VDD#163	XI1/net1#2	8.21861e-18
C1080	PHI#23	XI3/XI1/Q#2	2.86692e-17
C1081	SOUT0#8	VDD#173	7.25049e-18
C1082	GND#100	SOUT2#9	2.67289e-18
C1083	XI0/XI1/Q#9	XI0/XI1/XI4/net24#3	1.58103e-18
C1084	GND#62	SOUT2#18	3.58773e-18
C1085	XI2/XI1/Q#9	XI2/XI1/Q#3	2.18451e-18
C1086	XI3/XI1/D#20	VDD#109	2.76988e-18
C1087	SOUT0#5	CIN#4	4.20801e-18
C1088	net21#14	XI2/XI0/XI1/net2#2	1.85354e-18
C1089	XI1/XI1/XI4/net24#9	XI1/XI1/XI4/PHINOT#3	8.28164e-18
C1090	VDD#149	XI2/XI0/XI0/ANOT	2.05454e-18
C1091	VDD#148	net14#7	3.76854e-18
C1092	XI3/XI0/XI0/BNOT#5	SOUT3#1	4.41626e-18
C1093	PHI#11	XI1/XI1/XI4/net24	8.89281e-18
C1094	GND#96	net21#3	3.66677e-18
C1095	VDD#12	XI0/net1#2	1.29263e-17
C1096	RST#11	XI3/XI1/D#6	1.04408e-17
C1097	XI1/XI0/XI0/BNOT#11	net7#9	3.59305e-18
C1098	XI1/XI1/Q#5	VDD#40	6.36626e-17
C1099	VDD#26	SOUT0#22	3.78854e-17
C1100	GND#110	net7#3	3.66677e-18
C1101	XI2/XI1/Q#6	VDD#66	1.63056e-17
C1102	XI1/XI1/Q#7	VDD#124	1.95651e-18
C1103	VDD#123	VDD	4.74455e-17
C1104	GND#12	XI0/XI1/D	3.7665e-18
C1105	net21#19	VDD#94	1.37441e-17
C1106	CIN#9	SOUT0#9	3.7545e-17
C1107	GND#120	XI3/XI0/XI1/net2	2.76367e-18
C1108	VDD#160	VDD	2.30186e-17
C1109	XI0/XI1/D#6	XI0/XI1/D#5	4.49187e-18
C1110	XI3/XI1/D#4	VDD#109	2.24036e-18
C1111	XI0/XI0/XI0/BNOT#10	SOUT0#2	7.16694e-18
C1112	net21#8	XI3/XI0/XI0/BNOT#14	8.83203e-18
C1113	XI3/XI1/XI4/PHINOT#2	XI3/XI1/XI4/net24	3.28269e-17
C1114	XI2/XI1/XI4/PHINOT#9	PHI#15	1.27134e-18
C1115	RST#2	GND#152	4.18468e-18
C1116	XI3/XI0/XI0/BNOT#5	XI3/XI0/XI0/BNOT#6	8.47836e-18
C1117	VDD#171	XI0/XI0/XI0/ANOT	2.05454e-18
C1118	XI0/XI1/XI4/PHINOT#9	PHI#2	1.01564e-16
C1119	RST#9	XI2/net1#2	1.10422e-17
C1120	XI3/XI1/Q#12	XI3/XI1/XI4/net24#12	1.90043e-17
C1121	GND#36	XI1/XI0/XI0/ANOT#3	2.55369e-18
C1122	GND#129	SOUT2#16	1.37047e-17
C1123	GND#138	SOUT1#16	1.37047e-17
C1124	GND#38	XI1/XI1/XI4/net24#3	3.76841e-18
C1125	VDD#14	VDD#131	1.16687e-17
C1126	XI0/XI1/XI4/net24#2	XI0/XI1/Q#12	1.3891e-17
C1127	GND#119	VDD#134	1.10177e-17
C1128	XI2/net1#4	XI2/XI0/XI1/net2#3	1.41355e-18
C1129	GND#94	XI3/XI0/XI0/ANOT#3	4.34667e-18
C1130	XI0/XI1/D#14	GND#151	6.94823e-18
C1131	RST#2	GND#151	6.31281e-18
C1132	XI1/XI0/XI0/ANOT#6	SOUT1#3	2.75761e-18
C1133	XI0/XI0/XI0/BNOT#4	VDD#169	2.37247e-18
C1134	VDD#133	RST#13	1.68597e-17
C1135	XI1/XI1/XI4/net24#11	VDD	4.65294e-18
C1136	GND#46	net14#3	3.96405e-18
C1137	GND#74	XI3/XI1/D#14	2.68363e-17
C1138	SOUT3#11	XI3/net1#16	1.59072e-18
C1139	XI2/XI1/Q#7	XI2/XI1/XI4/net24	6.2497e-18
C1140	GND#132	XI2/XI1/XI4/net24#6	1.96676e-17
C1141	XI0/XI1/Q#7	XI0/XI1/Q#6	6.45394e-18
C1142	GND#131	XI2/XI1/D#2	5.80251e-18
C1143	XI0/net1#9	CIN#8	1.55592e-17
C1144	SOUT1#20	GND#137	1.26093e-17
C1145	XI1/net1#9	VDD	1.98755e-17
C1146	XI3/XI1/D#2	XI3/XI1/XI4/net24#2	4.04498e-17
C1147	VDD#34	SOUT1#1	4.22292e-18
C1148	XI1/net1#4	VDD	2.62325e-17
C1149	net7#19	VDD#34	6.27963e-18
C1150	XI1/XI1/XI4/net24#12	XI1/XI1/Q#2	2.89847e-18
C1151	VDD#80	net21	5.53658e-18
C1152	GND#66	SOUT2#9	5.27208e-18
C1153	GND#93	net21#9	4.17672e-18
C1154	XI1/XI0/XI0/BNOT#14	XI1/XI0/XI0/BNOT#4	7.00366e-18
C1155	VDD#52	SOUT1#22	3.78854e-17
C1156	VDD#76	XI2/XI0/XI1/net2#2	8.46721e-18
C1157	XI0/XI1/XI4/net24#9	XI0/XI1/XI4/net24#13	6.59037e-18
C1158	SOUT2#20	RST#8	1.76518e-17
C1159	SOUT2#16	SOUT2#18	1.30402e-17
C1160	VDD#64	XI2/net1#2	1.29263e-17
C1161	SOUT2#24	XI2/XI0/XI0/ANOT#3	2.93467e-18
C1162	VDD#162	VDD#38	1.0238e-17
C1163	net21#21	VDD#147	6.72863e-18
C1164	SOUT3#6	net21#5	3.39838e-18
C1165	GND#46	XI2/XI0/XI0/ANOT#6	4.05316e-17
C1166	GND#60	XI2/XI1/Q#9	3.30192e-17
C1167	GND#68	net21#3	3.96405e-18
C1168	SOUT3#4	net21#4	4.68557e-18
C1169	COUT#7	GND#119	1.4419e-17
C1170	XI1/XI1/Q#11	XI1/XI1/XI4/net24#12	2.96161e-17
C1171	VDD#155	RST#8	2.35653e-17
C1172	XI3/XI0/XI0/BNOT#4	VDD#136	2.37247e-18
C1173	XI1/XI1/XI4/net24#6	XI1/XI1/XI4/PHINOT#3	5.17189e-18
C1174	GND#66	GND#99	8.15798e-18
C1175	XI0/XI1/D#19	GND#149	1.63017e-18
C1176	PHI#5	XI0/XI1/Q#2	2.73644e-17
C1177	GND#113	VDD#167	1.84065e-17
C1178	GND#18	SOUT0#18	3.58773e-18
C1179	VDD#52	VDD#51	1.35961e-17
C1180	XI2/XI0/XI1/net2#15	SOUT2#20	5.36179e-18
C1181	XI1/XI0/XI1/net2#15	SOUT1#20	5.36179e-18
C1182	XI1/net1#4	VDD#160	1.4412e-17
C1183	SOUT1#4	net7#4	4.68557e-18
C1184	VDD#42	VDD#161	1.0979e-17
C1185	net7#15	XI0/XI0/XI1/net2#2	3.27874e-18
C1186	net21	SOUT3#1	3.65393e-18
C1187	VDD#170	VDD#169	1.8229e-17
C1188	SOUT3#16	SOUT3#18	1.30402e-17
C1189	RST#5	net7#4	1.53357e-17
C1190	XI2/XI1/Q#11	XI2/XI1/XI4/net24#12	2.96161e-17
C1191	VDD#68	XI2/net1#9	2.69821e-18
C1192	XI0/XI1/D#4	VDD#130	2.24036e-18
C1193	XI1/XI1/XI4/net24#9	XI1/XI1/D#17	7.89635e-18
C1194	COUT#7	VDD#136	6.72863e-18
C1195	SOUT2#3	XI2/XI0/XI0/BNOT#2	1.91621e-18
C1196	XI0/XI1/D#15	RST#2	4.36037e-17
C1197	XI2/XI1/Q#5	XI2/XI1/XI4/net24	3.34152e-18
C1198	SOUT2#16	XI2/XI1/Q#3	4.25775e-18
C1199	GND#24	net7#3	3.96405e-18
C1200	VDD#74	XI2/XI1/Q	4.68876e-18
C1201	XI0/XI1/D#17	XI0/XI1/Q#11	1.88867e-17
C1202	net21#17	XI3/net1#2	4.32779e-17
C1203	VDD#175	CIN#13	3.06108e-18
C1204	XI3/XI1/XI4/PHINOT#4	VDD#111	1.16528e-17
C1205	XI3/XI1/Q#9	XI3/XI1/XI4/net24#3	1.58103e-18
C1206	RST#11	net21#4	1.53357e-17
C1207	XI2/net1#4	VDD#149	1.4412e-17
C1208	XI3/XI1/D#19	XI3/XI1/XI4/net24#9	4.55106e-18
C1209	GND#64	XI2/XI0/XI1/net2	4.49691e-18
C1210	net21#15	RST#11	4.68358e-17
C1211	GND#131	XI2/XI1/D	2.42413e-18
C1212	GND#80	XI3/XI0/XI0/ANOT#3	2.55369e-18
C1213	GND#140	XI1/XI1/D#17	1.58396e-18
C1214	GND#88	GND#92	8.15798e-18
C1215	VDD#36	XI1/net1#2	1.39754e-17
C1216	XI2/XI1/D#14	GND#54	1.28303e-17
C1217	SOUT1#18	XI1/XI1/Q#2	5.04785e-18
C1218	XI3/XI1/Q#6	XI3/XI1/XI4/net24	1.04447e-18
C1219	RST#11	GND#125	1.95518e-17
C1220	VDD#122	VDD	8.65204e-17
C1221	GND#115	XI0/net1#16	1.74589e-17
C1222	VDD#165	RST#6	4.10956e-18
C1223	XI3/XI1/D#2	XI3/XI1/XI4/PHINOT#3	3.94365e-17
C1224	GND#16	XI0/XI1/Q#9	3.30192e-17
C1225	XI0/XI1/Q#6	VDD#14	1.63056e-17
C1226	XI0/XI1/XI4/net24#11	XI0/XI1/Q	4.03173e-18
C1227	SOUT1#11	XI1/XI0/XI0/BNOT#14	3.25292e-18
C1228	VDD#159	VDD	2.13492e-17
C1229	XI1/XI1/D#2	XI1/XI1/XI4/PHINOT#3	3.94365e-17
C1230	SOUT1#11	XI1/net1#16	1.59072e-18
C1231	XI2/XI1/Q#12	XI2/XI1/XI4/net24#13	1.81832e-17
C1232	RST#11	GND#76	1.18488e-17
C1233	XI2/XI1/XI4/net24#11	SOUT2#14	9.24112e-18
C1234	XI1/XI0/XI0/BNOT#7	XI1/XI0/XI0/BNOT#8	4.0203e-18
C1235	XI0/XI0/XI0/ANOT#4	VDD#8	2.2775e-17
C1236	XI2/XI1/XI4/PHINOT#2	PHI#14	2.96218e-17
C1237	RST#5	GND#20	1.13456e-17
C1238	VDD#145	VDD	4.3336e-17
C1239	XI1/XI0/XI0/ANOT#9	SOUT1#3	2.35212e-17
C1240	XI0/XI0/XI0/BNOT#14	SOUT0#22	8.52113e-18
C1241	XI0/XI1/XI4/net24#13	XI0/XI1/XI4/net24#2	1.71266e-17
C1242	VDD#66	XI2/XI1/XI4/PHINOT	3.64808e-18
C1243	SOUT2#11	XI2/XI0/XI0/BNOT#14	3.25292e-18
C1244	GND#24	XI1/XI0/XI0/ANOT#6	4.05316e-17
C1245	VDD#113	VDD	5.73405e-17
C1246	GND#123	GND#122	9.26445e-18
C1247	GND#117	CIN#3	3.66677e-18
C1248	net14#3	SOUT2#3	7.17245e-18
C1249	VDD#52	VDD	1.04322e-17
C1250	XI0/XI0/XI0/BNOT#7	SOUT0#3	5.63912e-18
C1251	VDD#94	SOUT3#7	8.24977e-18
C1252	VDD#142	net21#19	3.06108e-18
C1253	VDD#166	GND#144	1.78524e-17
C1254	VDD#115	XI2/XI1/Q	4.97335e-18
C1255	VDD#158	VDD	4.07404e-17
C1256	GND#141	XI1/XI1/XI4/net24#6	1.96676e-17
C1257	XI1/XI1/D#17	XI1/XI1/XI4/net24#12	8.08047e-18
C1258	VDD#176	RST#3	4.10956e-18
C1259	XI0/XI0/XI0/BNOT#5	SOUT0#2	1.8238e-17
C1260	net7	SOUT1#1	3.65393e-18
C1261	GND#52	XI2/XI1/D#14	2.68363e-17
C1262	XI3/XI1/Q#12	XI3/XI1/XI4/net24#13	1.81832e-17
C1263	SOUT0#8	SOUT0#11	8.1418e-18
C1264	net7#19	VDD#163	1.34565e-17
C1265	PHI#2	XI0/XI1/XI4/PHINOT#4	4.3751e-18
C1266	SOUT1#14	XI1/XI1/Q	7.83548e-18
C1267	XI1/XI1/XI4/net24#11	PHI#10	7.57347e-18
C1268	VDD#154	RST#9	4.10956e-18
C1269	SOUT1#14	VDD	8.86864e-18
C1270	XI1/net1#9	net7#8	1.55592e-17
C1271	XI0/XI1/XI4/net24	XI0/XI1/D#4	2.39789e-18
C1272	XI2/XI0/XI0/BNOT#5	SOUT2#1	4.41626e-18
C1273	GND#56	XI2/XI1/D#2	9.24969e-18
C1274	RST#2	XI0/net1#2	3.74826e-18
C1275	PHI#18	XI2/XI1/Q#3	3.05252e-18
C1276	VDD#52	VDD#158	1.09613e-17
C1277	SOUT0#8	XI0/XI0/XI0/ANOT	2.40961e-17
C1278	net14#10	VDD	8.95824e-18
C1279	GND#106	VDD#156	1.84065e-17
C1280	RST#5	XI1/net1#2	3.74826e-18
C1281	VDD#16	VDD#15	1.68878e-17
C1282	XI0/XI0/XI1/net2#15	net7#15	8.93527e-18
C1283	XI0/net1#4	VDD#170	1.37422e-18
C1284	SOUT0#24	XI0/XI0/XI0/BNOT#11	2.12646e-17
C1285	VDD#50	net14#10	5.51165e-17
C1286	SOUT0#20	net7#14	1.77949e-16
C1287	SOUT2#19	XI2/XI1/Q#3	5.30351e-18
C1288	SOUT0#22	GND#113	2.23064e-17
C1289	RST#12	XI3/net1#3	2.67237e-18
C1290	VDD#173	SOUT0#6	4.21273e-18
C1291	SOUT1#22	VDD	9.33159e-18
C1292	net14#12	SOUT1#20	2.00237e-17
C1293	VDD#117	XI2/XI1/XI4/PHINOT	4.411e-18
C1294	GND#56	XI2/XI1/D	3.7665e-18
C1295	SOUT1#20	VDD	7.57963e-18
C1296	SOUT2#10	net14#9	4.46078e-17
C1297	SOUT1#10	net7#9	4.46078e-17
C1298	XI3/XI1/XI4/net24#2	XI3/XI1/XI4/PHINOT#3	1.97764e-17
C1299	VDD#139	SOUT3#7	2.63522e-18
C1300	VDD#52	XI1/XI0/XI0/BNOT#3	8.47855e-18
C1301	VDD#159	XI1/XI0/XI1/net2#15	3.53013e-18
C1302	XI3/XI1/D#19	XI3/XI1/XI4/PHINOT#3	2.23795e-18
C1303	SOUT1#10	net7#8	3.40191e-18
C1304	VDD#169	XI0/XI0/XI1/net2#3	3.05777e-18
C1305	XI1/net1#4	VDD#50	8.38893e-18
C1306	COUT#1	XI3/XI0/XI1/net2#2	5.88268e-18
C1307	XI2/XI0/XI0/ANOT#4	VDD#60	2.2775e-17
C1308	net14#21	VDD	1.1147e-17
C1309	SOUT0#11	CIN#8	1.51494e-17
C1310	VDD#144	GND#126	1.78524e-17
C1311	XI2/XI1/XI4/net24#6	GND#56	3.31614e-17
C1312	VDD#60	XI2/XI0/XI0/BNOT#5	5.45774e-17
C1313	VDD#149	net14#6	4.16751e-18
C1314	XI1/XI1/XI4/net24#9	XI1/XI1/XI4/PHINOT#2	1.74823e-18
C1315	net14#14	VDD	1.10481e-17
C1316	net7#14	RST#5	4.02246e-17
C1317	XI3/XI1/D#17	XI3/XI1/XI4/PHINOT#3	8.962e-19
C1318	GND#139	PHI#12	5.83194e-18
C1319	SOUT3#11	XI3/net1#9	2.44574e-17
C1320	XI0/XI1/XI4/net24#11	SOUT0#14	9.24112e-18
C1321	XI1/XI0/XI0/BNOT#2	XI1/XI0/XI0/ANOT#2	6.90696e-17
C1322	SOUT1#16	SOUT1#17	4.09771e-18
C1323	GND#106	VDD	2.72001e-17
C1324	GND#138	SOUT1#18	1.34133e-17
C1325	GND#108	XI1/net1#16	1.74589e-17
C1326	GND#95	XI3/XI0/XI0/BNOT#7	1.31853e-17
C1327	GND#107	XI1/net1#16	9.27251e-18
C1328	XI1/XI1/XI4/net24#2	XI1/XI1/XI4/PHINOT#3	1.97764e-17
C1329	net7#19	SOUT1#2	6.17276e-17
C1330	VDD#94	XI3/net1#9	2.69821e-18
C1331	XI1/XI1/XI4/PHINOT#6	PHI#9	9.47309e-18
C1332	XI1/XI1/D#2	XI1/XI1/XI4/net24#4	1.54296e-18
C1333	XI3/XI1/XI4/net24#11	XI3/XI1/Q	4.03173e-18
C1334	GND#128	XI2/XI0/XI1/net2#2	1.86055e-18
C1335	SOUT0#14	SOUT0#15	6.95608e-18
C1336	RST#11	net21#12	7.49192e-18
C1337	XI0/XI0/XI0/BNOT#14	XI0/XI0/XI0/BNOT#4	7.00366e-18
C1338	VDD#105	GND#118	1.79196e-17
C1339	SOUT3#22	net21#8	5.05993e-18
C1340	XI2/XI1/D#14	XI2/net1	2.44048e-18
C1341	COUT#5	GND#119	1.08364e-16
C1342	VDD#155	VDD	7.78897e-17
C1343	XI1/XI1/Q#7	XI1/XI1/Q#5	9.68451e-18
C1344	VDD#141	XI3/net1#3	2.93418e-18
C1345	VDD#40	XI1/XI1/D#3	1.58831e-18
C1346	XI3/XI1/D#14	GND#124	6.94823e-18
C1347	XI0/net1#16	XI0/XI0/XI0/ANOT#2	2.38906e-18
C1348	SOUT3#18	VDD#105	2.18537e-17
C1349	VDD#50	XI1/XI0/XI1/net2#3	5.00211e-18
C1350	XI3/XI0/XI0/BNOT	XI3/XI0/XI0/ANOT#3	4.63673e-17
C1351	VDD#119	VDD	9.39951e-17
C1352	XI2/XI1/Q#6	VDD#117	4.14214e-18
C1353	GND#62	SOUT2#16	4.02471e-17
C1354	XI3/XI1/D#10	XI3/net1#2	7.8648e-18
C1355	PHI#17	XI2/XI1/Q	1.20146e-17
C1356	GND#129	SOUT2#19	3.10131e-18
C1357	PHI#5	XI0/XI1/XI4/net24	8.89281e-18
C1358	SOUT3#19	SOUT3#18	3.98821e-17
C1359	CIN#13	VDD#174	1.34565e-17
C1360	XI1/XI0/XI1/net2#2	SOUT1#20	1.29961e-17
C1361	RST#11	GND#123	9.12929e-18
C1362	GND#10	SOUT0#4	4.09574e-18
C1363	VDD#78	net14#7	4.04071e-18
C1364	XI0/XI0/XI0/BNOT#2	XI0/XI0/XI0/ANOT#3	9.13179e-18
C1365	VDD#54	VDD	1.49508e-17
C1366	GND#2	CIN#3	3.96405e-18
C1367	XI1/XI1/Q#12	XI1/XI1/XI4/PHINOT#2	2.90831e-18
C1368	net7#15	SOUT0#20	8.75531e-17
C1369	VDD#154	VDD	7.27918e-17
C1370	GND#76	SOUT3#4	4.09574e-18
C1371	VDD#112	XI2/XI1/Q#2	2.47832e-18
C1372	XI1/XI0/XI0/ANOT#9	net7#2	4.97779e-17
C1373	XI1/XI0/XI0/ANOT#6	XI1/XI0/XI0/BNOT#7	5.36256e-18
C1374	XI2/net1#2	SOUT2#5	3.43763e-18
C1375	XI1/XI1/Q#9	SOUT1#16	1.50594e-18
C1376	VDD#12	SOUT0#6	4.07255e-18
C1377	VDD#44	XI1/XI1/XI4/net24	1.58831e-18
C1378	XI0/XI1/Q#6	XI0/XI1/D#20	8.17481e-17
C1379	net7	SOUT1#2	2.69766e-18
C1380	net14	SOUT2#1	3.65393e-18
C1381	VDD#72	net14#6	4.0872e-18
C1382	SOUT3#2	VDD#140	3.04495e-18
C1383	XI3/XI1/XI4/net24#4	XI3/XI1/Q#12	2.8824e-17
C1384	XI1/XI1/XI4/net24#11	XI1/XI1/XI4/net24#10	7.53548e-18
C1385	net7#17	XI1/XI1/D#14	5.73862e-18
C1386	XI2/XI1/D#4	VDD#70	4.83878e-18
C1387	XI3/XI1/Q#9	PHI#24	4.56241e-18
C1388	SOUT2#19	SOUT2#18	3.98821e-17
C1389	RST#8	net14#4	1.53357e-17
C1390	XI1/XI0/XI0/BNOT	XI1/XI0/XI0/ANOT#3	4.63673e-17
C1391	VDD#88	XI3/net1#3	3.96888e-18
C1392	GND#122	XI3/XI1/D#2	5.80251e-18
C1393	VDD#56	VDD	1.68456e-17
C1394	XI2/XI0/XI0/BNOT#11	SOUT2#22	7.23396e-18
C1395	XI1/XI1/XI4/net24#4	XI1/XI1/Q#12	2.8824e-17
C1396	SOUT3#10	XI3/XI0/XI0/BNOT#11	3.84272e-17
C1397	XI0/XI1/Q#5	VDD#131	1.53345e-17
C1398	XI0/XI1/D#19	XI0/XI1/XI4/PHINOT#3	2.23795e-18
C1399	VDD#118	VDD	1.32558e-16
C1400	CIN#1	VDD	2.10514e-17
C1401	RST#6	XI1/net1#3	2.67237e-18
C1402	SOUT3#5	net21#5	4.43091e-17
C1403	net21#17	SOUT3#5	2.7909e-17
C1404	XI1/XI1/D#4	VDD#44	4.83878e-18
C1405	VDD#57	VDD	2.12045e-17
C1406	XI3/XI1/D#19	XI3/XI1/XI4/net24#6	1.52492e-17
C1407	GND#40	SOUT1#16	4.02471e-17
C1408	XI2/XI1/D#2	XI2/XI1/XI4/PHINOT#3	3.94365e-17
C1409	VDD#149	VDD#72	1.0238e-17
C1410	RST#3	VDD	2.21559e-17
C1411	XI1/XI1/Q#5	VDD#124	1.53345e-17
C1412	SOUT3#18	PHI#23	1.77809e-17
C1413	XI3/XI0/XI0/ANOT#6	XI3/XI0/XI0/BNOT#7	5.36256e-18
C1414	GND#10	GND#150	1.0238e-17
C1415	GND#138	SOUT1#19	3.10131e-18
C1416	XI2/XI1/D#19	XI2/XI1/XI4/PHINOT#2	8.83178e-18
C1417	PHI#1	VDD	2.39701e-17
C1418	XI1/XI1/D#19	PHI#9	2.62196e-18
C1419	SOUT0#2	VDD#174	4.81645e-18
C1420	SOUT0#1	VDD	7.47753e-18
C1421	VDD#14	VDD#18	3.93119e-17
C1422	SOUT3#10	net21#8	3.40191e-18
C1423	GND#86	GND#120	8.84679e-18
C1424	VDD#134	VDD	4.33201e-17
C1425	XI2/XI0/XI0/ANOT#4	VDD	9.31981e-18
C1426	GND#106	net14#21	1.0327e-16
C1427	XI0/net1#3	VDD	4.47542e-18
C1428	SOUT3#16	SOUT3#17	4.09771e-18
C1429	SOUT1#18	GND#137	3.44305e-17
C1430	VDD#106	VDD	5.73743e-17
C1431	VDD#143	RST#12	4.10956e-18
C1432	XI3/XI1/D	XI3/XI1/XI4/net24#3	2.52567e-18
C1433	XI0/XI1/Q#9	PHI#6	4.56241e-18
C1434	COUT#6	XI3/XI0/XI1/net2#2	3.27874e-18
C1435	XI2/net1#16	SOUT2#24	5.33627e-17
C1436	SOUT0#6	VDD	1.22001e-17
C1437	SOUT1#5	RST#5	3.79452e-17
C1438	GND#134	GND#48	9.24934e-18
C1439	XI3/XI1/Q#7	XI3/XI1/Q#5	9.68451e-18
C1440	VDD#150	XI2/net1#9	1.70357e-18
C1441	net7#12	SOUT0#16	2.93637e-18
C1442	XI1/XI1/XI4/PHINOT#9	PHI#9	1.27134e-18
C1443	XI0/XI1/XI4/PHINOT	VDD	1.47213e-17
C1444	SOUT0#5	RST#2	3.79452e-17
C1445	VDD#154	VDD#57	1.02424e-17
C1446	GND#8	GND#7	7.83801e-18
C1447	XI2/net1#4	XI2/XI0/XI1/net2#15	3.27011e-17
C1448	net14#12	SOUT1#16	2.93637e-18
C1449	XI0/XI1/XI4/net24	VDD	9.38808e-18
C1450	GND#95	SOUT3#3	5.38904e-18
C1451	RST#7	XI2/net1	3.14306e-18
C1452	net7#19	SOUT1#8	2.94542e-17
C1453	VDD#72	XI2/net1#4	3.90041e-17
C1454	XI2/net1#16	XI2/XI0/XI0/BNOT#11	1.66841e-17
C1455	PHI#8	VDD#30	6.00445e-18
C1456	VDD#94	XI3/XI0/XI0/ANOT	4.13602e-18
C1457	RST#5	GND#139	6.19589e-18
C1458	XI2/XI1/XI4/PHINOT#9	VDD	4.78049e-18
C1459	net14#2	VDD#54	3.99391e-18
C1460	XI3/XI0/XI0/BNOT#5	VDD#141	1.54612e-17
C1461	CIN#11	RST#2	7.73029e-18
C1462	SOUT0#18	XI0/XI1/Q#2	5.04785e-18
C1463	VDD#149	XI2/XI0/XI1/net2#15	1.7071e-18
C1464	VDD#70	XI2/XI1/D#3	6.45552e-18
C1465	SOUT0#7	VDD	3.25902e-18
C1466	XI0/XI1/D#2	XI0/XI1/XI4/net24#3	1.40726e-18
C1467	COUT#5	RST#13	4.02246e-17
C1468	XI0/XI0/XI0/BNOT#14	CIN#7	1.32694e-17
C1469	net7#8	XI1/XI0/XI0/BNOT#4	3.19507e-18
C1470	XI0/XI1/Q#6	XI0/XI1/XI4/net24	1.04447e-18
C1471	XI2/XI1/D#17	XI2/XI1/Q#12	5.03747e-17
C1472	RST#11	GND#129	7.91186e-18
C1473	XI2/XI1/XI4/PHINOT#4	VDD	2.14306e-17
C1474	SOUT1#24	XI1/XI0/XI0/BNOT#2	5.12165e-17
C1475	SOUT0#18	XI0/XI1/Q#3	1.55626e-18
C1476	XI0/XI0/XI0/ANOT#4	XI0/XI0/XI0/BNOT#5	1.1098e-17
C1477	XI0/XI0/XI0/ANOT	VDD	5.29805e-18
C1478	GND#123	SOUT3#4	3.19662e-18
C1479	XI1/XI0/XI0/BNOT#11	SOUT1#22	7.23396e-18
C1480	XI2/XI1/D#10	VDD	1.26139e-17
C1481	CIN#6	VDD	1.13782e-17
C1482	VDD#144	XI2/XI0/XI1/net2#2	1.25381e-18
C1483	XI0/XI1/XI4/PHINOT#6	XI0/XI1/D#19	8.37816e-18
C1484	VDD#98	XI3/XI0/XI1/net2#3	1.01229e-18
C1485	net14#9	SOUT2#9	3.7545e-17
C1486	XI0/XI1/D#3	VDD	4.65131e-18
C1487	CIN#1	SOUT0#2	2.69766e-18
C1488	XI3/XI1/Q#11	PHI#24	1.32498e-17
C1489	VDD#151	VDD#64	1.0238e-17
C1490	GND#150	SOUT0#4	3.19662e-18
C1491	PHI#4	VDD	5.74562e-18
C1492	XI1/XI1/XI4/net24#2	XI1/XI1/XI4/net24#4	1.52005e-18
C1493	XI3/XI1/D#15	XI3/net1#2	3.59645e-18
C1494	VDD#171	CIN#6	4.16751e-18
C1495	XI3/XI1/XI4/net24#6	XI3/XI1/XI4/net24#5	6.84508e-18
C1496	VDD#164	net7#19	3.06108e-18
C1497	CIN#7	VDD	5.19162e-18
C1498	SOUT0#24	XI0/XI0/XI0/ANOT#2	7.14175e-18
C1499	PHI#11	XI1/XI1/XI4/PHINOT#2	4.78246e-17
C1500	XI0/XI1/Q	VDD	2.04814e-17
C1501	VDD#46	XI1/net1#4	3.90041e-17
C1502	SOUT2#20	GND#128	1.26093e-17
C1503	SOUT2#11	net14#8	1.51116e-17
C1504	XI0/XI0/XI0/BNOT#2	XI0/XI0/XI0/ANOT#2	6.90696e-17
C1505	SOUT0#24	XI0/XI0/XI0/ANOT#3	2.93467e-18
C1506	RST#2	GND#147	7.22408e-18
C1507	VDD#153	VDD	1.8633e-17
C1508	VDD#104	VDD#136	1.09613e-17
C1509	GND#141	XI1/XI1/D#19	1.45214e-17
C1510	VDD#160	XI1/XI0/XI1/net2#15	1.7071e-18
C1511	XI0/XI0/XI0/BNOT#3	VDD	4.09757e-18
C1512	XI0/XI1/D#2	XI0/XI1/XI4/net24#4	1.54296e-18
C1513	VDD#96	XI3/XI1/XI4/net24#11	6.32412e-17
C1514	GND#141	XI1/XI1/D#2	3.24657e-18
C1515	XI1/XI1/D	XI1/XI1/XI4/net24#3	2.52567e-18
C1516	VDD#8	SOUT0#1	4.22292e-18
C1517	XI1/XI0/XI1/net2#16	SOUT1#5	2.87586e-18
C1518	VDD#139	XI3/XI0/XI0/ANOT	1.82797e-18
C1519	XI0/XI0/XI1/net2#3	VDD	8.39596e-18
C1520	VDD#66	XI2/XI1/XI4/net24	6.41722e-18
C1521	GND#64	net21#12	4.0234e-17
C1522	GND#56	GND#60	1.79944e-17
C1523	XI2/XI0/XI0/BNOT#4	net14#7	2.43471e-17
C1524	XI1/XI1/XI4/net24#6	XI1/XI1/D	1.8988e-18
C1525	GND#93	SOUT3#9	2.67289e-18
C1526	VDD#102	COUT#1	5.51165e-17
C1527	VDD#133	COUT#5	1.42169e-18
C1528	net7	VDD	2.10514e-17
C1529	XI0/XI1/D#20	VDD#18	2.68757e-17
C1530	RST#9	XI2/net1#3	2.67237e-18
C1531	SOUT1#10	SOUT1#22	5.91301e-18
C1532	XI1/XI1/Q#7	XI1/XI1/XI4/PHINOT	1.21362e-17
C1533	XI2/XI1/XI4/net24#2	XI2/XI1/XI4/PHINOT#3	1.97764e-17
C1534	XI1/XI1/XI4/net24#6	XI1/XI1/D#17	1.49998e-18
C1535	VDD#116	XI2/XI1/D#3	4.10481e-18
C1536	XI2/XI0/XI0/ANOT#9	SOUT2#2	2.69483e-18
C1537	RST#6	VDD	2.21559e-17
C1538	net14#10	net14#11	7.3184e-18
C1539	VDD#139	XI3/net1#9	1.70357e-18
C1540	VDD#148	SOUT2#20	2.94846e-18
C1541	SOUT2#14	PHI#17	1.23563e-17
C1542	XI3/XI1/XI4/net24	XI3/XI1/D#4	2.39789e-18
C1543	XI0/XI1/D#19	GND#151	3.09843e-17
C1544	XI1/XI1/Q#6	XI1/XI1/XI4/PHINOT#2	2.75539e-18
C1545	PHI#7	VDD	2.39701e-17
C1546	XI1/XI0/XI1/net2#16	net7#5	2.63779e-17
C1547	XI0/XI1/XI4/net24#11	XI0/XI1/XI4/net24#10	7.53548e-18
C1548	XI2/XI0/XI0/BNOT#5	VDD	8.81368e-18
C1549	XI2/XI1/D#4	VDD#116	2.24036e-18
C1550	GND#78	XI3/XI1/D#2	9.24969e-18
C1551	VDD#20	XI0/XI0/XI1/net2#16	1.4293e-18
C1552	COUT#1	SOUT3#20	4.66076e-17
C1553	SOUT1#1	VDD	7.47753e-18
C1554	RST#13	GND#120	1.51603e-17
C1555	net7#2	XI1/XI0/XI0/ANOT#4	3.09365e-18
C1556	SOUT3#14	SOUT3#18	1.77557e-17
C1557	XI3/XI1/XI4/net24#4	XI3/XI1/Q#11	1.49839e-17
C1558	VDD#152	VDD	1.94359e-17
C1559	XI1/net1#3	VDD	4.47542e-18
C1560	XI3/net1#16	XI3/XI0/XI0/ANOT#2	2.38906e-18
C1561	XI2/XI1/D#14	GND#133	6.94823e-18
C1562	PHI#23	VDD#100	5.40385e-18
C1563	XI3/XI0/XI0/BNOT#14	net21#7	1.32694e-17
C1564	XI2/XI0/XI0/ANOT#2	XI2/XI0/XI0/BNOT#10	7.01434e-17
C1565	XI0/XI1/D#19	XI0/XI1/XI4/PHINOT#2	8.83178e-18
C1566	XI2/XI0/XI1/net2#16	SOUT2#6	5.16806e-18
C1567	SOUT1#6	VDD	1.22001e-17
C1568	XI3/XI1/D#14	SOUT3#5	7.88532e-18
C1569	XI1/XI0/XI1/net2#13	RST#5	2.21589e-17
C1570	XI1/XI1/D#17	XI1/XI1/Q#12	5.03747e-17
C1571	GND#147	XI0/XI1/Q#3	2.16945e-18
C1572	GND#30	XI1/net1	4.05515e-18
C1573	GND#72	SOUT3#3	4.36955e-18
C1574	XI0/XI1/D#2	XI0/XI1/D#17	3.60142e-18
C1575	SOUT1#11	XI1/net1#9	2.44574e-17
C1576	GND#72	XI3/XI0/XI0/BNOT#7	4.05316e-17
C1577	XI2/XI1/D#17	PHI#18	1.97458e-18
C1578	XI1/XI1/XI4/PHINOT	VDD	1.47213e-17
C1579	GND#120	SOUT3#18	1.34133e-17
C1580	GND#114	GND#22	9.65661e-18
C1581	XI0/XI1/Q#11	PHI#6	1.32498e-17
C1582	net21#8	XI3/XI0/XI0/BNOT#4	3.19507e-18
C1583	VDD#2	XI0/XI0/XI0/ANOT#4	5.51165e-17
C1584	XI1/XI1/XI4/net24	VDD	9.38808e-18
C1585	CIN#2	SOUT0#3	2.27501e-18
C1586	XI2/net1#9	XI2/XI0/XI0/ANOT	1.29015e-18
C1587	XI3/XI1/D#19	GND#124	3.09843e-17
C1588	SOUT3#5	net21#4	4.20801e-18
C1589	net14#19	VDD	7.38122e-18
C1590	XI2/XI0/XI0/BNOT#11	net14#8	1.64202e-18
C1591	VDD#159	XI1/XI0/XI1/net2#2	4.26212e-18
C1592	XI0/XI1/XI4/net24#9	XI0/XI1/D#17	7.89635e-18
C1593	XI2/XI0/XI0/BNOT#10	SOUT2#2	7.16694e-18
C1594	SOUT1#7	VDD	3.25902e-18
C1595	XI1/XI1/D#4	VDD#123	2.24036e-18
C1596	VDD#20	CIN#6	4.0872e-18
C1597	XI1/XI1/XI4/PHINOT#4	XI1/XI1/XI4/PHINOT#5	5.34824e-18
C1598	net14#17	VDD	6.33291e-18
C1599	XI1/XI1/D#20	VDD#44	2.68757e-17
C1600	XI3/XI0/XI1/net2#16	net21#5	2.63779e-17
C1601	VDD#22	SOUT0#14	5.47763e-17
C1602	XI1/XI0/XI0/ANOT	VDD	5.29805e-18
C1603	SOUT3#8	XI3/XI0/XI0/ANOT	2.40961e-17
C1604	SOUT0#8	VDD#16	1.33308e-17
C1605	XI0/XI0/XI0/BNOT#2	XI0/XI0/XI0/BNOT#9	1.3821e-17
C1606	VDD#117	XI2/XI1/XI4/net24	4.3074e-18
C1607	net7#6	VDD	1.13782e-17
C1608	XI1/XI1/D#20	XI1/XI1/XI4/net24#12	1.97297e-17
C1609	PHI#23	XI3/XI1/XI4/net24	8.89281e-18
C1610	VDD#152	VDD#62	1.0238e-17
C1611	XI0/XI1/D#19	GND#12	2.48425e-18
C1612	XI1/XI1/D#3	VDD	4.65131e-18
C1613	XI0/XI0/XI0/ANOT#6	SOUT0#3	2.75761e-18
C1614	RST#8	GND#52	1.03647e-17
C1615	XI3/XI1/D#15	XI3/net1	1.96101e-17
C1616	VDD#46	XI1/XI0/XI1/net2#16	1.4293e-18
C1617	GND#143	GND#26	9.24934e-18
C1618	VDD#151	VDD	2.56909e-17
C1619	PHI#10	VDD	5.74562e-18
C1620	XI0/XI1/D#17	XI0/XI1/XI4/net24#12	8.08047e-18
C1621	XI1/XI1/Q#5	XI1/XI1/XI4/PHINOT	8.79316e-18
C1622	VDD#165	VDD#31	1.02424e-17
C1623	XI1/XI0/XI0/BNOT#5	SOUT1#1	4.41626e-18
C1624	GND#34	GND#38	1.79944e-17
C1625	RST#5	GND#32	1.18488e-17
C1626	net7#7	VDD	5.19162e-18
C1627	XI0/XI0/XI0/BNOT#5	VDD#174	1.54612e-17
C1628	VDD#140	XI3/net1#2	9.35443e-18
C1629	VDD#171	VDD#20	1.0238e-17
C1630	XI2/XI1/XI4/net24#4	XI2/XI1/Q#12	2.8824e-17
C1631	VDD#20	XI0/XI0/XI1/net2#3	1.01229e-18
C1632	GND#88	SOUT3#9	5.27208e-18
C1633	XI1/XI1/Q	VDD	2.04814e-17
C1634	XI0/XI1/XI4/PHINOT#3	XI0/XI1/D	3.80638e-17
C1635	SOUT2#20	RST#11	2.00652e-17
C1636	GND#86	XI3/XI0/XI1/net2	4.49691e-18
C1637	XI1/XI0/XI0/BNOT#3	VDD	4.09757e-18
C1638	VDD#68	VDD#150	1.0979e-17
C1639	XI0/XI1/Q#6	VDD#131	4.14214e-18
C1640	XI1/XI1/D#10	XI1/net1#2	7.8648e-18
C1641	GND#30	GND#142	1.02095e-17
C1642	SOUT1#11	net7#8	1.51116e-17
C1643	XI0/XI0/XI1/net2#13	XI0/XI0/XI1/net2	2.66668e-18
C1644	XI1/XI0/XI1/net2#3	VDD	8.39596e-18
C1645	VDD#16	SOUT0#7	8.24977e-18
C1646	XI0/XI0/XI1/net2#13	CIN#4	2.31785e-18
C1647	XI0/XI1/XI4/net24#6	XI0/XI1/XI4/net24#5	6.84508e-18
C1648	net7#17	VDD#163	2.19992e-17
C1649	VDD#119	PHI#14	2.63987e-17
C1650	XI1/XI0/XI0/ANOT#4	net7	6.05749e-18
C1651	RST#6	XI1/net1#2	1.10422e-17
C1652	GND#130	net14#4	3.80483e-18
C1653	XI0/XI1/D#17	XI0/XI1/XI4/net24#4	3.52091e-17
C1654	VDD#4	XI0/XI1/XI4/PHINOT#4	5.55471e-17
C1655	net14	VDD	2.10514e-17
C1656	XI0/XI1/XI4/net24#4	XI0/XI1/Q#11	1.49839e-17
C1657	XI0/net1#16	SOUT0#24	5.33627e-17
C1658	net7#10	XI0/XI0/XI1/net2#3	6.65581e-18
C1659	GND#76	GND#123	1.0238e-17
C1660	SOUT1#5	net7#4	4.20801e-18
C1661	VDD#152	XI2/net1#3	2.93418e-18
C1662	RST#9	VDD	2.21559e-17
C1663	GND#130	GND#60	1.0238e-17
C1664	RST#8	GND#135	1.64699e-17
C1665	XI0/XI1/Q#9	XI0/XI1/Q#11	1.53602e-18
C1666	XI0/XI1/D#14	RST#2	5.02859e-17
C1667	net21#10	SOUT2#20	4.66076e-17
C1668	XI2/XI1/Q#7	VDD	1.11747e-17
C1669	PHI#13	VDD	2.39701e-17
C1670	XI1/XI0/XI0/BNOT#10	net7#2	2.58085e-18
C1671	SOUT2#14	SOUT2#18	1.77557e-17
C1672	GND#40	SOUT1#18	3.58773e-18
C1673	XI1/XI1/XI4/net24#13	XI1/XI1/XI4/PHINOT#2	2.64065e-17
C1674	GND#131	XI2/XI1/D#17	1.58396e-18
C1675	XI2/net1#16	SOUT2#10	4.33498e-18
C1676	XI2/XI1/Q#5	VDD	1.57977e-17
C1677	GND#116	XI0/XI0/XI0/BNOT#7	1.08055e-17
C1678	SOUT2#1	VDD	7.47753e-18
C1679	GND#121	GND#82	1.0238e-17
C1680	XI3/XI0/XI0/BNOT#7	XI3/XI0/XI0/ANOT#9	4.40775e-18
C1681	GND#146	RST#5	2.41904e-17
C1682	XI2/XI0/XI0/BNOT#9	SOUT2#22	1.14498e-17
C1683	XI2/net1#3	VDD	4.47542e-18
C1684	XI2/XI0/XI0/ANOT#4	net14	6.05749e-18
C1685	XI2/XI1/D#17	XI2/XI1/Q#9	7.82323e-18
C1686	SOUT2#6	VDD	1.22001e-17
C1687	VDD#92	VDD#110	1.16687e-17
C1688	XI0/XI1/XI4/PHINOT	XI0/XI1/XI4/net24	7.48941e-17
C1689	XI3/XI1/Q#9	XI3/XI1/Q#8	3.3441e-18
C1690	XI2/XI0/XI0/ANOT#2	net14#8	2.9337e-18
C1691	XI2/net1#4	XI2/XI0/XI1/net2#2	9.28475e-19
C1692	XI0/XI0/XI1/net2#13	net7#15	8.86742e-18
C1693	SOUT0#11	XI0/XI0/XI0/ANOT#2	1.22267e-18
C1694	XI0/XI0/XI0/BNOT#11	XI0/XI0/XI0/BNOT#9	1.98917e-17
C1695	XI0/net1#4	XI0/XI0/XI1/net2#15	3.27011e-17
C1696	XI2/XI1/XI4/PHINOT	VDD	1.47213e-17
C1697	XI0/XI0/XI1/net2#13	GND#148	1.3169e-17
C1698	SOUT0#10	CIN#8	3.40191e-18
C1699	VDD#92	XI3/XI1/D#3	1.58831e-18
C1700	XI0/net1#16	XI0/XI0/XI0/BNOT#11	1.66841e-17
C1701	GND#142	XI1/net1	4.15538e-18
C1702	XI3/XI1/D#17	XI3/XI1/Q#9	7.82323e-18
C1703	VDD#170	XI0/XI0/XI1/net2#15	3.53013e-18
C1704	XI2/XI1/XI4/net24	VDD	9.38808e-18
C1705	XI1/XI1/XI4/net24#9	XI1/XI1/D#2	3.0624e-17
C1706	XI2/XI1/XI4/PHINOT#6	XI2/XI1/D#19	8.37816e-18
C1707	GND#18	XI0/XI1/Q#3	4.41398e-18
C1708	XI0/XI0/XI0/BNOT#5	XI0/XI0/XI0/BNOT#6	8.47836e-18
C1709	XI3/XI1/XI4/net24#12	XI3/XI1/XI4/net24#4	1.1037e-18
C1710	SOUT1#18	XI1/XI1/Q#3	1.55626e-18
C1711	XI0/XI0/XI1/net2#2	SOUT0#20	1.29961e-17
C1712	XI2/XI0/XI0/ANOT#4	SOUT2#2	5.09768e-18
C1713	XI0/XI1/XI4/net24#2	XI0/XI1/XI4/net24#4	1.52005e-18
C1714	GND#149	XI0/XI1/D#2	5.80251e-18
C1715	SOUT2#7	VDD	3.25902e-18
C1716	XI0/net1#4	VDD#24	8.38893e-18
C1717	XI3/XI0/XI1/net2#15	COUT#1	6.82353e-18
C1718	GND#100	SOUT2#10	7.13064e-18
C1719	VDD#117	VDD	8.4118e-17
C1720	XI3/XI0/XI0/BNOT#10	net21#2	2.58085e-18
C1721	XI2/XI0/XI0/ANOT	VDD	5.29805e-18
C1722	XI3/XI1/Q#7	XI3/XI1/Q#6	6.45394e-18
C1723	PHI#5	XI0/XI1/XI4/PHINOT#2	4.78246e-17
C1724	XI2/XI0/XI0/BNOT#11	net14#9	3.59305e-18
C1725	VDD#30	XI1/XI1/XI4/PHINOT#4	5.55471e-17
C1726	SOUT0#24	XI0/XI0/XI0/BNOT#9	6.98011e-18
C1727	GND#123	XI3/XI1/XI4/PHINOT#3	3.59673e-18
C1728	XI0/XI1/XI4/net24#11	VDD#22	1.81691e-17
C1729	VDD#34	XI1/XI0/XI0/BNOT#5	5.45774e-17
C1730	net14#6	VDD	1.13782e-17
C1731	XI0/XI1/D#14	GND#10	1.28303e-17
C1732	SOUT3#16	XI3/XI1/Q#3	4.25775e-18
C1733	GND#6	CIN#3	1.73249e-18
C1734	VDD#158	XI1/XI0/XI1/net2#3	3.05777e-18
C1735	XI2/XI1/XI4/net24#9	XI2/XI1/XI4/net24#13	6.59037e-18
C1736	XI2/net1#2	SOUT2#6	1.96305e-17
C1737	GND#114	XI0/net1#16	9.27251e-18
C1738	XI1/XI0/XI0/BNOT#11	XI1/XI0/XI0/BNOT#9	1.98917e-17
C1739	XI2/XI1/D#3	VDD	4.65131e-18
C1740	XI0/XI1/XI4/net24#6	GND#12	3.31614e-17
C1741	VDD#62	XI2/net1#3	3.96888e-18
C1742	XI0/XI0/XI0/ANOT#4	CIN#1	6.05749e-18
C1743	PHI#16	VDD	5.74562e-18
C1744	VDD#172	SOUT0#7	2.63522e-18
C1745	SOUT2#11	XI2/net1#16	1.59072e-18
C1746	VDD#150	VDD	1.44935e-17
C1747	XI0/XI0/XI0/ANOT#9	CIN#2	4.9727e-17
C1748	XI3/XI1/XI4/net24#11	VDD#109	1.56401e-17
C1749	net14#7	VDD	5.19162e-18
C1750	XI1/XI1/Q#9	SOUT1#19	5.37314e-18
C1751	XI2/XI0/XI0/BNOT#9	net14#8	9.80156e-17
C1752	XI3/net1#9	VDD#137	7.01142e-18
C1753	XI2/XI1/D#19	XI2/XI1/D#2	1.57987e-18
C1754	XI2/XI1/D#19	GND#131	1.63017e-18
C1755	VDD#170	XI0/XI0/XI1/net2#2	4.26212e-18
C1756	XI2/XI1/Q	VDD	2.04814e-17
C1757	XI0/XI0/XI0/ANOT#9	SOUT0#3	2.35212e-17
C1758	COUT#6	SOUT3#20	8.75531e-17
C1759	XI2/XI1/Q#6	VDD	9.99629e-18
C1760	XI2/XI0/XI0/BNOT#5	SOUT2#2	1.8238e-17
C1761	XI1/XI1/XI4/net24#11	VDD#48	1.81691e-17
C1762	XI2/net1#9	VDD#148	7.01142e-18
C1763	XI2/net1#16	XI2/XI0/XI0/BNOT#9	1.54391e-17
C1764	PHI#20	VDD#82	6.00445e-18
C1765	XI2/XI0/XI0/BNOT#3	VDD	4.09757e-18
C1766	VDD#50	XI1/XI0/XI1/net2#2	8.46721e-18
C1767	XI2/XI1/XI4/net24#11	XI2/XI1/XI4/net24#10	7.53548e-18
C1768	VDD#18	XI0/XI1/D#3	6.45552e-18
C1769	XI2/XI0/XI1/net2#3	VDD	8.39596e-18
C1770	XI2/XI0/XI1/net2#16	VDD	3.04753e-18
C1771	net21	VDD	2.10514e-17
C1772	XI1/XI0/XI0/BNOT#7	XI1/XI0/XI0/ANOT#9	4.40775e-18
C1773	XI3/XI0/XI1/net2#13	net21#4	2.31785e-18
C1774	GND#84	SOUT3#18	3.58773e-18
C1775	GND#146	VDD#167	1.10177e-17
C1776	RST#12	VDD	2.21559e-17
C1777	XI2/XI1/Q#12	XI2/XI1/D#20	2.28141e-17
C1778	RST#8	GND#133	6.31281e-18
C1779	VDD#90	XI3/net1#2	1.29263e-17
C1780	GND#99	net21#21	1.0327e-16
C1781	RST#5	XI0/XI0/XI1/net2	1.51821e-17
C1782	XI0/XI1/Q#9	SOUT0#16	1.50594e-18
C1783	RST#3	XI0/net1#2	1.10422e-17
C1784	SOUT2#18	GND#128	3.44305e-17
C1785	XI3/XI1/XI4/PHINOT	XI3/XI1/XI4/net24	7.48941e-17
C1786	VDD#126	GND#144	2.2414e-17
C1787	PHI#19	VDD	2.39701e-17
C1788	SOUT0#8	VDD#172	5.47184e-18
C1789	net14#21	GND#137	1.4419e-17
C1790	VDD#57	RST#9	5.42714e-18
C1791	SOUT2#16	SOUT2#19	1.38255e-17
C1792	net7#12	SOUT0#20	2.00237e-17
C1793	net7#15	XI0/XI0/XI1/net2	7.48119e-18
C1794	XI2/XI1/D#20	VDD	3.67809e-18
C1795	VDD#126	XI0/XI1/Q	2.29584e-18
C1796	XI2/XI1/Q#9	XI2/XI1/Q#8	3.3441e-18
C1797	SOUT3#1	VDD	7.47753e-18
C1798	VDD#66	VDD#117	1.16687e-17
C1799	VDD#31	RST#6	5.42714e-18
C1800	XI0/net1#9	XI0/XI0/XI0/ANOT	1.29015e-18
C1801	GND#140	GND#34	1.01892e-17
C1802	SOUT3#24	XI3/XI0/XI0/BNOT#2	5.12165e-17
C1803	XI3/net1#3	VDD	4.47542e-18
C1804	GND#108	XI1/XI0/XI0/BNOT#2	3.63595e-18
C1805	XI1/XI1/D#4	PHI#10	1.07136e-17
C1806	RST#5	GND#141	9.12929e-18
C1807	XI2/XI0/XI1/net2#16	net14#5	2.63779e-17
C1808	SOUT3#6	VDD	1.22001e-17
C1809	XI0/XI1/Q#6	PHI#5	4.16718e-17
C1810	XI1/XI1/XI4/PHINOT#2	PHI#8	2.96218e-17
C1811	XI1/XI1/Q#9	XI1/XI1/XI4/net24#3	1.58103e-18
C1812	XI3/XI1/XI4/PHINOT	VDD	1.47213e-17
C1813	GND#132	XI2/XI1/D#19	1.45214e-17
C1814	VDD#76	SOUT2#20	4.21807e-18
C1815	SOUT1#20	VDD#158	2.36869e-17
C1816	VDD#112	GND#126	2.2414e-17
C1817	XI3/XI1/XI4/net24	VDD	9.38808e-18
C1818	XI2/XI1/Q#7	XI2/XI1/Q#6	6.45394e-18
C1819	SOUT3#18	XI3/XI1/Q#2	5.04785e-18
C1820	XI2/XI1/XI4/PHINOT#4	XI2/XI1/XI4/PHINOT#5	5.34824e-18
C1821	XI1/XI1/D#15	XI1/net1#2	3.59645e-18
C1822	GND#8	GND#151	1.02095e-17
C1823	XI0/XI1/XI4/net24#13	PHI#5	9.76906e-18
C1824	SOUT3#19	XI3/XI1/Q#3	5.30351e-18
C1825	XI3/XI1/XI4/net24#9	XI3/XI1/XI4/PHINOT#3	8.28164e-18
C1826	CIN#11	VDD#174	2.19992e-17
C1827	net21#17	XI3/XI1/D#14	5.73862e-18
C1828	SOUT3#7	VDD	3.25902e-18
C1829	XI1/XI0/XI0/BNOT#9	SOUT1#22	1.14498e-17
C1830	XI0/XI1/XI4/PHINOT#6	PHI#3	9.47309e-18
C1831	XI3/XI1/D#6	RST#10	5.54809e-18
C1832	XI3/XI1/Q#9	XI3/XI1/Q#3	2.18451e-18
C1833	XI3/XI0/XI0/ANOT	VDD	5.29805e-18
C1834	XI3/XI0/XI0/ANOT#4	net21	6.05749e-18
C1835	XI1/XI1/XI4/net24#9	XI1/XI1/Q#12	4.7443e-18
C1836	VDD#116	PHI#16	4.96959e-18
C1837	XI0/XI0/XI0/BNOT#11	CIN#8	1.64202e-18
C1838	XI0/XI1/XI4/net24#12	XI0/XI1/XI4/net24#4	1.1037e-18
C1839	GND#84	XI3/XI1/Q#2	5.13993e-18
C1840	net21#6	VDD	1.13782e-17
C1841	XI0/XI1/XI4/PHINOT#2	PHI#2	2.96218e-17
C1842	XI3/XI0/XI0/BNOT#2	XI3/XI0/XI0/ANOT#3	9.13179e-18
C1843	VDD#116	VDD	4.74455e-17
C1844	XI1/XI1/Q#7	XI1/XI1/XI4/PHINOT#2	9.18965e-19
C1845	SOUT2#5	net14#4	4.20801e-18
C1846	XI3/XI1/D#3	VDD	4.65131e-18
C1847	XI2/XI0/XI1/net2#15	XI2/XI0/XI1/net2#2	6.41939e-18
C1848	XI3/XI0/XI0/ANOT#9	net21#2	4.97779e-17
C1849	VDD#130	XI0/XI1/D#3	4.10481e-18
C1850	VDD#149	VDD	2.30186e-17
C1851	XI3/XI0/XI0/ANOT#3	net21#9	1.57734e-18
C1852	PHI#22	VDD	5.74562e-18
C1853	XI3/XI0/XI0/BNOT#2	XI3/XI0/XI0/ANOT#2	6.90696e-17
C1854	net7#19	XI1/XI0/XI0/ANOT#2	1.52499e-17
C1855	SOUT3#20	RST#13	3.33183e-17
C1856	XI3/XI0/XI0/ANOT#2	XI3/XI0/XI0/BNOT#10	7.01434e-17
C1857	GND#102	SOUT2#3	5.38904e-18
C1858	VDD#166	RST#5	2.35653e-17
C1859	GND#149	GND#12	1.01892e-17
C1860	XI3/XI1/D#2	XI3/XI1/XI4/net24#4	1.54296e-18
C1861	GND#10	GND#9	7.9864e-18
C1862	GND#14	XI0/XI0/XI0/ANOT#2	4.32997e-18
C1863	net21#7	VDD	5.19162e-18
C1864	SOUT1	XI1/XI1/Q	2.71859e-18
C1865	net14#14	XI1/XI0/XI1/net2#2	1.85354e-18
C1866	GND#66	SOUT2#10	1.12163e-17
C1867	SOUT0	XI0/XI1/Q	2.71859e-18
C1868	XI3/XI0/XI0/BNOT#7	XI3/XI0/XI0/BNOT#8	4.0203e-18
C1869	XI3/XI1/Q	VDD	2.04814e-17
C1870	SOUT2#24	XI2/XI0/XI0/BNOT#2	5.12165e-17
C1871	SOUT1#11	XI1/XI0/XI0/ANOT	8.09714e-18
C1872	XI3/XI0/XI0/BNOT#3	VDD	4.09757e-18
C1873	XI3/XI0/XI1/net2#2	SOUT3#20	1.29961e-17
C1874	GND#134	XI2/XI1/XI4/PHINOT#6	1.36671e-17
C1875	XI1/net1#16	XI1/XI0/XI0/ANOT#2	2.38906e-18
C1876	GND#137	VDD#156	1.10177e-17
C1877	XI1/XI1/XI4/net24#6	XI1/XI1/D#2	9.87705e-18
C1878	SOUT0#6	CIN#6	3.8605e-18
C1879	SOUT0#20	VDD#169	2.36869e-17
C1880	SOUT1#22	XI1/XI0/XI0/BNOT#4	3.05405e-18
C1881	CIN#8	XI0/XI0/XI0/BNOT#4	3.19507e-18
C1882	XI2/XI1/D#19	GND#133	3.09843e-17
C1883	XI3/XI0/XI1/net2#3	VDD	8.39596e-18
C1884	XI2/XI0/XI0/BNOT#9	net14#19	1.54043e-17
C1885	XI1/XI0/XI0/BNOT#5	VDD#163	1.54612e-17
C1886	SOUT2	XI2/XI1/Q	2.71859e-18
C1887	GND#110	GND#24	8.47392e-18
C1888	GND#42	GND#138	8.84679e-18
C1889	GND#22	GND#21	7.74457e-18
C1890	VDD#175	VDD#174	1.68962e-17
C1891	XI0/XI1/XI4/net24#9	XI0/XI1/Q#12	4.7443e-18
C1892	XI2/XI1/XI4/net24#11	VDD	4.65294e-18
C1893	net7#17	XI1/net1#2	4.32779e-17
C1894	VDD#148	VDD#147	1.8229e-17
C1895	GND#12	XI0/XI1/D#2	9.24969e-18
C1896	XI0/XI0/XI1/net2#15	SOUT0#5	5.93898e-18
C1897	net21#2	SOUT3#2	1.06752e-17
C1898	XI0/XI1/XI4/PHINOT#4	XI0/XI1/XI4/PHINOT#5	5.34824e-18
C1899	VDD#83	RST#12	5.42714e-18
C1900	GND#92	COUT	9.09265e-18
C1901	VDD#147	XI2/XI0/XI1/net2#2	1.54384e-18
C1902	net14#8	XI2/XI0/XI0/BNOT#14	8.83203e-18
C1903	VDD#174	XI0/net1#2	8.21861e-18
C1904	XI2/XI1/Q#6	VDD#116	1.9494e-18
C1905	XI3/XI0/XI0/BNOT#14	XI3/XI0/XI0/BNOT#4	7.00366e-18
C1906	XI2/XI1/D#6	RST#7	5.54809e-18
C1907	GND#115	XI0/XI0/XI0/BNOT	2.7139e-18
C1908	XI2/net1#9	VDD	1.98755e-17
C1909	XI1/XI1/D#19	XI1/XI1/XI4/net24#9	4.55106e-18
C1910	SOUT3#6	net21#6	3.8605e-18
C1911	GND#116	GND#6	8.36698e-18
C1912	SOUT2#14	XI2/XI1/Q	7.83548e-18
C1913	SOUT0#4	CIN#4	4.68557e-18
C1914	VDD#175	XI0/XI1/D#10	1.29802e-17
C1915	net14#15	XI1/XI0/XI1/net2	7.48119e-18
C1916	XI2/net1#4	VDD	2.62325e-17
C1917	RST#2	XI0/net1	2.28596e-17
C1918	VDD#96	XI3/XI1/XI4/net24	1.58831e-18
C1919	VDD#78	XI2/XI0/XI0/BNOT#3	8.47855e-18
C1920	net7#12	XI0/XI0/XI1/net2	5.18165e-18
C1921	XI1/XI1/Q#7	XI1/XI1/XI4/net24	6.2497e-18
C1922	SOUT2#2	VDD#152	4.81645e-18
C1923	GND#99	VDD#145	1.84065e-17
C1924	VDD#5	RST#3	5.42714e-18
C1925	GND#119	VDD#133	7.65081e-17
C1926	VDD#44	XI1/XI1/XI4/net24#11	6.32412e-17
C1927	SOUT3	XI3/XI1/Q	2.71859e-18
C1928	XI0/XI1/D#10	CIN#11	1.25206e-17
C1929	XI3/XI0/XI1/net2#15	COUT#6	8.93527e-18
C1930	PHI#2	VDD#4	6.00445e-18
C1931	XI3/net1#4	XI3/XI0/XI1/net2#3	1.41355e-18
C1932	XI3/XI1/D#17	XI3/XI1/Q#11	1.88867e-17
C1933	XI3/XI1/XI4/net24#6	XI3/XI1/XI4/PHINOT#3	5.17189e-18
C1934	VDD#24	XI0/XI0/XI1/net2#2	8.46721e-18
C1935	VDD#76	XI2/XI0/XI1/net2#3	5.00211e-18
C1936	XI2/XI0/XI0/BNOT#10	net14#19	1.41727e-16
C1937	VDD#66	XI2/XI1/XI4/net24#13	1.09794e-18
C1938	SOUT3#10	SOUT3#22	5.91301e-18
C1939	XI1/XI1/XI4/net24#6	XI1/XI1/XI4/net24#5	6.84508e-18
C1940	XI3/XI0/XI0/BNOT#10	XI3/XI0/XI0/ANOT#9	7.21709e-17
C1941	CIN#2	XI0/XI0/XI0/ANOT#4	3.09365e-18
C1942	net21#15	SOUT2#20	8.75531e-17
C1943	XI3/XI1/XI4/net24#6	GND#78	3.31614e-17
C1944	SOUT2#19	XI2/XI1/Q#2	6.59904e-18
C1945	XI3/XI1/D#2	XI3/XI1/XI4/net24#3	1.40726e-18
C1946	SOUT0#10	SOUT0#22	5.91301e-18
C1947	VDD#44	VDD#123	1.16687e-17
C1948	XI2/net1#4	net14#6	1.35025e-17
C1949	GND#101	XI2/XI0/XI0/BNOT	2.7139e-18
C1950	XI1/XI0/XI0/BNOT#11	net7#8	1.64202e-18
C1951	XI1/XI0/XI0/ANOT#6	GND#28	1.48844e-17
C1952	XI1/XI1/Q#12	XI1/XI1/D#20	2.28141e-17
C1953	GND#130	XI2/XI1/XI4/net24#3	4.14351e-18
C1954	XI2/net1#16	XI2/XI0/XI0/ANOT#2	2.38906e-18
C1955	COUT#3	SOUT3#20	2.00237e-17
C1956	XI2/XI0/XI0/BNOT#14	SOUT2#22	8.52113e-18
C1957	XI3/net1#4	VDD#137	1.37422e-18
C1958	XI3/XI1/XI4/net24#3	PHI#24	4.68747e-17
C1959	GND#20	net7#12	4.0234e-17
C1960	GND#150	XI0/XI1/XI4/PHINOT#3	3.59673e-18
C1961	VDD#153	VDD#152	1.68962e-17
C1962	XI3/XI1/D#19	XI3/XI1/XI4/PHINOT#2	8.83178e-18
C1963	VDD#141	VDD#88	1.0238e-17
C1964	VDD#137	net21#7	3.76854e-18
C1965	XI1/XI1/D#20	VDD#123	2.76988e-18
C1966	COUT#7	VDD#134	7.44569e-18
C1967	XI0/XI1/XI4/PHINOT#9	PHI#3	1.27134e-18
C1968	VDD#56	PHI#13	6.76392e-18
C1969	VDD#170	SOUT0#20	2.94846e-18
C1970	GND#50	SOUT2#3	4.36955e-18
C1971	GND#36	XI1/XI0/XI0/BNOT#2	1.48416e-18
C1972	XI1/XI0/XI0/BNOT#2	XI1/XI0/XI0/ANOT#3	9.13179e-18
C1973	SOUT1#10	XI1/XI0/XI0/BNOT#4	2.61929e-18
C1974	XI1/XI0/XI0/BNOT#9	net7#19	1.54043e-17
C1975	XI1/XI1/D#20	XI1/XI1/XI4/net24#11	1.30924e-17
C1976	XI0/XI1/D#20	VDD#130	2.76988e-18
C1977	XI1/net1#2	SOUT1#5	3.43763e-18
C1978	XI1/XI1/XI4/net24#11	XI1/XI1/Q	4.03173e-18
C1979	XI3/XI1/XI4/net24#9	XI3/XI1/D#17	7.89635e-18
C1980	XI2/XI1/D#17	XI2/XI1/Q#11	1.88867e-17
C1981	XI2/XI0/XI0/ANOT#6	XI2/XI0/XI0/BNOT#7	5.36256e-18
C1982	VDD#115	VDD	8.65204e-17
C1983	XI3/XI1/Q#6	PHI#23	4.16718e-17
C1984	XI2/XI1/D#10	net14#17	1.25206e-17
C1985	XI3/XI1/Q#11	PHI#23	1.16343e-17
C1986	XI1/XI0/XI1/net2#13	XI1/XI0/XI1/net2	2.66668e-18
C1987	VDD#148	VDD	2.13492e-17
C1988	XI1/XI1/Q#5	XI1/XI1/XI4/net24	3.34152e-18
C1989	GND#138	XI1/XI1/Q#3	2.16945e-18
C1990	net21#2	XI3/XI0/XI0/ANOT#4	3.09365e-18
C1991	GND#146	VDD#166	7.65081e-17
C1992	XI2/XI1/D#4	PHI#17	2.70764e-17
C1993	SOUT3#24	XI3/XI0/XI0/BNOT#11	2.12646e-17
C1994	SOUT0#20	XI0/XI0/XI1/net2#3	1.51276e-18
C1995	SOUT3#10	XI3/XI0/XI0/BNOT#4	2.61929e-18
C1996	XI3/XI1/XI4/net24#2	XI3/XI1/XI4/net24#4	1.52005e-18
C1997	PHI#5	XI0/XI1/Q#7	3.39064e-17
C1998	CIN#11	XI0/XI1/D#14	5.73862e-18
C1999	XI1/XI0/XI0/ANOT#9	net7#19	6.99675e-18
C2000	XI1/XI1/XI4/net24#9	XI1/XI1/XI4/net24#13	6.59037e-18
C2001	XI1/XI0/XI1/net2#16	XI1/net1#4	3.40431e-17
C2002	PHI#23	XI3/XI1/XI4/PHINOT#2	4.78246e-17
C2003	SOUT0#14	VDD#129	1.16528e-17
C2004	XI0/XI1/D#17	XI0/XI1/XI4/net24#2	6.90619e-18
C2005	XI3/XI0/XI0/BNOT#2	XI3/XI0/XI0/BNOT#9	1.3821e-17
C2006	XI1/XI0/XI0/ANOT#3	net7#9	1.57734e-18
C2007	XI1/XI1/Q#12	XI1/XI1/XI4/net24#12	1.90043e-17
C2008	SOUT1#8	SOUT1#11	8.1418e-18
C2009	XI0/XI0/XI0/BNOT#9	CIN#8	9.80977e-17
C2010	XI2/XI1/XI4/net24#11	XI2/XI1/D#3	3.27281e-18
C2011	SOUT3#7	XI3/XI0/XI0/ANOT	5.39732e-17
C2012	GND#34	XI1/XI1/XI4/PHINOT#3	2.02958e-18
C2013	XI2/XI1/Q#6	XI2/XI1/XI4/net24	1.04447e-18
C2014	VDD#30	PHI#7	6.76392e-18
C2015	XI0/XI1/D#19	XI0/XI1/D#2	1.57987e-18
C2016	XI0/net1#2	SOUT0#5	3.43763e-18
C2017	net14#10	XI1/XI0/XI1/net2#3	6.65581e-18
C2018	VDD#82	PHI#19	6.76392e-18
C2019	XI2/XI1/D#2	XI2/XI1/XI4/PHINOT#2	1.00039e-18
C2020	XI0/XI1/Q#12	XI0/XI1/XI4/net24#12	1.90043e-17
C2021	net14#12	XI1/XI0/XI1/net2	5.18165e-18
C2022	VDD#78	VDD	1.04322e-17
C2023	VDD#40	XI1/XI1/XI4/PHINOT	3.64808e-18
C2024	XI1/XI1/D#19	GND#140	1.63017e-18
C2025	XI0/XI1/XI4/net24#6	XI0/XI1/D#17	1.49998e-18
C2026	SOUT2#11	XI2/net1#9	2.44574e-17
C2027	XI2/net1#4	VDD#148	1.37422e-18
C2028	VDD#36	net7#17	2.54235e-17
C2029	XI2/XI0/XI0/ANOT#9	net14#19	6.99675e-18
C2030	XI2/XI1/XI4/PHINOT#9	PHI#14	1.01564e-16
C2031	VDD#147	VDD	4.07404e-17
C2032	SOUT1#2	VDD#162	3.04495e-18
C2033	XI2/net1#9	XI2/XI0/XI0/BNOT#9	3.86468e-18
C2034	net7#12	GND#147	1.3363e-17
C2035	GND#14	XI0/XI0/XI0/BNOT	4.9463e-18
C2036	RST#11	GND#126	1.64699e-17
C2037	net21#21	GND#128	1.4419e-17
C2038	SOUT2#18	XI2/XI1/Q#3	1.55626e-18
C2039	XI2/XI1/XI4/net24#4	XI2/XI1/Q#11	1.49839e-17
C2040	XI0/XI1/D#20	XI0/XI1/XI4/net24#12	1.97297e-17
C2041	GND#58	XI2/XI0/XI0/BNOT	4.9463e-18
C2042	XI0/XI0/XI0/ANOT#4	VDD#176	1.1119e-17
C2043	GND#60	XI2/XI1/XI4/net24#3	3.76841e-18
C2044	VDD#100	XI3/XI1/Q	4.68876e-18
C2045	SOUT0#7	XI0/XI0/XI0/ANOT	5.39732e-17
C2046	SOUT2#14	VDD	8.86864e-18
C2047	XI2/XI1/D#19	GND#56	2.48425e-18
C2048	VDD#147	net21#10	1.49363e-17
C2049	XI2/XI1/D#15	XI2/net1	1.96101e-17
C2050	XI3/XI1/XI4/net24#11	XI3/XI1/D#4	3.45102e-18
C2051	SOUT1#14	PHI#11	1.23563e-17
C2052	net21#10	VDD	8.95824e-18
C2053	GND#114	CIN#9	4.17672e-18
C2054	XI3/net1#4	net21#5	1.24619e-17
C2055	XI2/XI1/Q#9	GND#62	1.37107e-17
C2056	XI2/XI1/Q#6	XI2/XI1/D#20	8.17481e-17
C2057	GND#100	SOUT2#22	9.0763e-18
C2058	XI1/XI1/D#2	XI1/XI1/XI4/net24#3	1.40726e-18
C2059	XI1/XI1/D#14	XI1/net1	2.44048e-18
C2060	VDD#140	SOUT3#6	4.21273e-18
C2061	XI2/XI1/D#19	XI2/XI1/XI4/PHINOT#3	2.23795e-18
C2062	XI1/XI1/XI4/net24#4	XI1/XI1/Q#11	1.49839e-17
C2063	VDD#42	VDD#41	1.68878e-17
C2064	GND#64	SOUT2#20	5.19922e-18
C2065	XI1/XI1/XI4/PHINOT	XI1/XI1/XI4/net24	7.48941e-17
C2066	XI1/XI1/XI4/net24#9	XI1/XI1/XI4/net24#2	7.14446e-18
C2067	RST#11	XI2/XI0/XI1/net2	1.51821e-17
C2068	XI3/XI1/XI4/net24	XI3/XI1/D#3	2.28624e-18
C2069	VDD#16	VDD#172	1.0979e-17
C2070	XI0/XI0/XI1/net2#13	SOUT0#5	2.17512e-17
C2071	SOUT2#22	VDD	9.33159e-18
C2072	SOUT0#11	XI0/net1#16	1.59072e-18
C2073	XI1/XI1/Q#11	SOUT1#19	7.03151e-18
C2074	VDD#22	SOUT0	4.09262e-18
C2075	VDD#10	XI0/net1#2	1.39754e-17
C2076	XI0/XI1/XI4/net24#9	XI0/XI1/XI4/PHINOT#3	8.28164e-18
C2077	COUT#3	COUT#4	4.31453e-18
C2078	VDD#16	XI0/XI0/XI0/ANOT	4.13602e-18
C2079	SOUT2#20	VDD	7.57963e-18
C2080	SOUT0	VDD#129	3.91522e-17
C2081	net21#14	RST#11	4.02246e-17
C2082	VDD#170	CIN#7	3.76854e-18
C2083	XI1/XI1/D#6	RST#4	5.54809e-18
C2084	XI0/XI0/XI0/BNOT#5	SOUT0#1	4.41626e-18
C2085	VDD#163	XI1/net1#3	2.93418e-18
C2086	XI2/XI1/Q#12	XI2/XI1/XI4/PHINOT#2	2.90831e-18
C2087	XI3/XI0/XI0/BNOT#7	SOUT3#3	5.63912e-18
C2088	RST#2	SOUT0#4	2.05565e-17
C2089	XI0/net1#9	VDD#171	3.67621e-17
C2090	net21#21	VDD	1.1147e-17
C2091	XI1/XI1/XI4/net24#6	GND#34	3.31614e-17
C2092	net14#17	RST#8	7.73029e-18
C2093	XI1/XI0/XI0/BNOT#9	net7#8	9.80156e-17
C2094	GND#149	XI0/XI1/D#17	1.58396e-18
C2095	VDD#159	VDD#158	1.8229e-17
C2096	SOUT0#20	GND#146	1.26093e-17
C2097	GND#54	SOUT2#4	4.09574e-18
C2098	XI3/XI1/D#17	XI3/XI1/XI4/net24#4	3.52091e-17
C2099	VDD#124	XI1/XI1/XI4/PHINOT	4.411e-18
C2100	VDD#108	XI3/XI1/Q	4.97335e-18
C2101	net21#14	VDD	1.10481e-17
C2102	GND#30	GND#29	7.83801e-18
C2103	VDD#68	SOUT2#7	8.24977e-18
C2104	XI1/XI1/XI4/PHINOT#4	VDD#125	1.16528e-17
C2105	XI2/XI1/XI4/PHINOT	XI2/XI1/XI4/net24	7.48941e-17
C2106	GND#76	GND#75	7.9864e-18
C2107	XI1/XI1/XI4/net24#2	XI1/XI1/Q#12	1.3891e-17
C2108	GND#40	XI1/XI1/Q#3	4.41398e-18
C2109	GND#99	VDD	2.72001e-17
C2110	XI0/XI1/XI4/PHINOT#4	VDD#132	1.16528e-17
C2111	XI0/XI0/XI1/net2#13	net7#12	3.2914e-18
C2112	XI3/XI0/XI1/net2#13	COUT#6	8.86742e-18
C2113	SOUT0#14	PHI#5	1.23563e-17
C2114	net14#14	GND#137	1.08364e-16
C2115	XI2/XI1/D#19	XI2/XI1/XI4/net24#9	4.55106e-18
C2116	VDD#66	VDD#70	3.93119e-17
C2117	GND#96	GND#68	8.47392e-18
C2118	SOUT3#22	XI3/XI0/XI0/BNOT#4	3.05678e-18
C2119	SOUT1#18	VDD#119	2.18537e-17
C2120	XI0/net1#16	XI0/XI0/XI0/BNOT#9	1.54391e-17
C2121	XI2/XI0/XI0/BNOT#2	XI2/XI0/XI0/ANOT#3	9.13179e-18
C2122	VDD#144	VDD	7.78897e-17
C2123	XI1/XI1/XI4/net24#3	PHI#12	4.68747e-17
C2124	XI3/XI1/XI4/net24#12	PHI#23	4.06087e-17
C2125	XI2/XI1/D#16	RST#8	5.13284e-17
C2126	VDD#54	XI2/XI0/XI0/ANOT#4	5.51165e-17
C2127	GND#6	XI0/XI0/XI0/BNOT#7	4.05316e-17
C2128	SOUT0#14	SOUT0	3.64962e-17
C2129	VDD#90	SOUT3#6	4.07255e-18
C2130	VDD#112	VDD	9.39951e-17
C2131	GND#86	COUT#3	4.0234e-17
C2132	XI0/net1#4	CIN#5	1.24619e-17
C2133	net7#12	net7#13	4.31453e-18
C2134	VDD#26	VDD#25	1.35961e-17
C2135	XI0/net1#4	XI0/XI0/XI1/net2#2	9.28475e-19
C2136	XI1/net1#4	XI1/XI0/XI1/net2#2	9.28475e-19
C2137	XI0/XI1/XI4/net24	XI0/XI1/D#3	2.28624e-18
C2138	XI3/XI1/D#17	XI3/XI1/XI4/net24#12	8.08047e-18
C2139	net21#15	XI2/XI0/XI1/net2	7.48119e-18
C2140	XI0/XI1/D#19	PHI#3	2.62196e-18
C2141	VDD#137	XI3/XI0/XI1/net2#15	3.53013e-18
C2142	RST#8	XI1/XI0/XI1/net2	1.51821e-17
C2143	VDD#137	SOUT3#20	2.94846e-18
C2144	SOUT1#8	VDD#162	7.25049e-18
C2145	XI2/XI1/XI4/net24#9	XI2/XI1/D#17	7.89635e-18
C2146	net7#2	VDD#28	3.99391e-18
C2147	VDD#80	VDD	1.49508e-17
C2148	XI1/net1#4	XI1/XI0/XI1/net2#15	3.27011e-17
C2149	GND#100	GND#66	9.65661e-18
C2150	XI3/net1#4	VDD#102	8.38893e-18
C2151	XI3/XI1/XI4/net24#6	XI3/XI1/D	1.8988e-18
C2152	net14#5	XI2/XI0/XI1/net2#2	4.87283e-18
C2153	XI1/net1#16	XI1/XI0/XI0/BNOT#11	1.66841e-17
C2154	SOUT3#8	SOUT3#11	8.1418e-18
C2155	XI1/XI0/XI0/BNOT#14	SOUT1#22	8.52113e-18
C2156	net7#17	VDD#162	6.83507e-18
C2157	XI3/XI1/Q#9	XI3/XI1/Q#11	1.53602e-18
C2158	VDD#143	VDD	7.27918e-17
C2159	XI1/XI1/Q#9	PHI#12	4.56241e-18
C2160	XI1/XI0/XI0/BNOT#10	XI1/XI0/XI0/ANOT#9	7.21709e-17
C2161	XI0/XI0/XI0/BNOT	XI0/XI0/XI0/ANOT#3	4.63673e-17
C2162	XI1/net1#16	SOUT1#10	4.33498e-18
C2163	XI3/net1#4	XI3/XI0/XI1/net2#15	3.27011e-17
C2164	SOUT0#20	XI0/XI0/XI1/net2	2.16801e-17
C2165	GND#130	XI2/XI1/D#17	4.75796e-18
C2166	XI1/XI1/XI4/PHINOT#6	XI1/XI1/D#19	8.37816e-18
C2167	VDD#173	VDD#12	1.0238e-17
C2168	SOUT3#11	XI3/XI0/XI0/ANOT	8.09714e-18
C2169	XI3/XI0/XI0/ANOT#4	XI3/XI0/XI0/BNOT#10	2.24348e-18
C2170	XI3/XI1/D#6	GND#125	1.65584e-17
C2171	XI3/net1#16	XI3/XI0/XI0/BNOT#11	1.66841e-17
C2172	XI0/XI0/XI0/ANOT#6	XI0/XI0/XI0/BNOT#7	5.36256e-18
C2173	VDD#36	XI1/net1#3	3.96888e-18
C2174	VDD#74	SOUT2#14	5.47763e-17
C2175	GND#93	XI3/net1#16	9.27251e-18
C2176	VDD#172	XI0/XI0/XI0/ANOT	1.82797e-18
C2177	XI0/XI1/D#4	PHI#4	1.07136e-17
C2178	VDD#150	SOUT2#7	2.63522e-18
C2179	VDD#119	XI1/XI1/Q	2.29584e-18
C2180	SOUT0	VDD#126	1.57577e-17
C2181	XI2/XI1/XI4/PHINOT#2	XI2/XI1/XI4/net24#2	5.77081e-17
C2182	XI0/XI0/XI0/ANOT#2	XI0/XI0/XI0/BNOT#10	7.01434e-17
C2183	RST	GND#152	1.67283e-17
C2184	XI2/XI1/XI4/PHINOT#2	XI2/XI1/XI4/net24	3.28269e-17
C2185	net14#17	XI2/XI1/D#14	5.73862e-18
C2186	GND#22	CIN#9	2.55369e-18
C2187	XI1/XI0/XI0/BNOT#2	XI1/XI0/XI0/BNOT#9	1.3821e-17
C2188	GND#96	XI3/XI0/XI0/ANOT#6	1.31853e-17
C2189	RST#11	XI3/net1#2	3.74826e-18
C2190	VDD#119	XI1/XI1/Q#2	2.47832e-18
C2191	CIN#13	SOUT0#2	6.17276e-17
C2192	PHI#14	XI2/XI1/XI4/PHINOT#4	4.3751e-18
C2193	GND#137	XI1/XI0/XI1/net2#2	1.86055e-18
C2194	CIN#8	XI0/XI0/XI0/BNOT#14	8.83203e-18
C2195	GND#48	XI2/XI1/XI4/PHINOT#6	4.0951e-17
C2196	XI3/XI1/D#19	XI3/XI1/D#2	1.57987e-18
C2197	net21#12	SOUT2#20	2.00237e-17
C2198	VDD#82	VDD	1.68456e-17
C2199	VDD#4	PHI#1	6.76392e-18
C2200	XI3/XI0/XI1/net2#13	GND#121	1.3169e-17
C2201	XI2/XI1/D#15	RST#8	4.36037e-17
C2202	net14#19	SOUT2#8	2.94542e-17
C2203	XI2/XI1/XI4/net24#12	XI2/XI1/XI4/net24#4	1.1037e-18
C2204	XI3/XI1/XI4/net24#6	XI3/XI1/D#17	1.49998e-18
C2205	VDD#111	VDD	1.32558e-16
C2206	SOUT1#24	XI1/XI0/XI0/ANOT#2	7.14175e-18
C2207	XI3/XI0/XI0/BNOT#10	net21#19	1.41727e-16
C2208	XI3/XI0/XI1/net2#15	net21#5	7.43893e-18
C2209	XI3/XI0/XI0/ANOT#6	net21#3	5.33566e-18
C2210	XI0/XI1/Q#9	SOUT0#19	5.37314e-18
C2211	VDD#83	VDD	2.12045e-17
C2212	net7#3	SOUT1#3	7.17245e-18
C2213	PHI#25	VDD	4.1237e-17
C2214	PHI#11	XI1/XI1/Q	1.20146e-17
C2215	XI0/net1#16	SOUT0#10	4.33498e-18
C2216	XI0/XI1/Q#5	XI0/XI1/Q#4	9.30041e-18
C2217	GND#148	CIN#4	3.80483e-18
C2218	SOUT3#24	XI3/XI0/XI0/BNOT#9	6.98011e-18
C2219	GND#132	SOUT2#4	3.19662e-18
C2220	XI0/XI1/XI4/net24#6	XI0/XI1/XI4/PHINOT#3	5.17189e-18
C2221	XI0/XI1/D#17	XI0/XI1/XI4/PHINOT#3	8.962e-19
C2222	XI0/XI1/D#6	GND#152	1.65584e-17
C2223	XI2/XI1/D#2	XI2/XI1/XI4/net24#3	1.40726e-18
C2224	net14#15	RST#8	4.68358e-17
C2225	COUT#6	RST#13	4.68358e-17
C2226	GND#108	GND#36	9.66245e-18
C2227	XI3/XI1/Q#9	SOUT3#16	1.50594e-18
C2228	VDD#152	XI2/net1#2	8.21861e-18
C2229	XI3/XI0/XI0/ANOT#4	VDD	9.31981e-18
C2230	GND#130	PHI#18	5.83194e-18
C2231	XI0/XI0/XI0/BNOT#10	CIN#2	2.58085e-18
C2232	XI2/XI1/XI4/net24#9	XI2/XI1/XI4/PHINOT#2	1.74823e-18
C2233	VDD#48	SOUT1	4.09262e-18
C2234	SOUT3#24	XI3/XI0/XI0/ANOT#2	7.14175e-18
C2235	GND#101	XI2/XI0/XI0/ANOT#3	4.34667e-18
C2236	XI1/XI0/XI0/BNOT#14	net7#7	1.32694e-17
C2237	VDD#104	net21#7	4.04071e-18
C2238	XI2/XI0/XI0/BNOT#5	net14#19	4.10074e-17
C2239	GND#64	GND#129	8.84679e-18
C2240	net7#14	XI0/XI0/XI1/net2#2	1.85354e-18
C2241	SOUT1	VDD#122	3.80499e-17
C2242	GND#117	XI0/XI0/XI0/ANOT#6	1.31853e-17
C2243	PHI#24	XI3/XI1/Q#3	3.05252e-18
C2244	SOUT1#6	net7#6	3.8605e-18
C2245	XI1/XI1/XI4/net24#12	XI1/XI1/XI4/net24#4	1.1037e-18
C2246	VDD#147	XI2/XI0/XI1/net2#3	3.05777e-18
C2247	XI2/XI1/Q#6	XI2/XI1/XI4/PHINOT#2	2.75539e-18
C2248	SOUT2#6	net14#6	3.8605e-18
C2249	net21#12	XI2/XI0/XI1/net2	5.18165e-18
C2250	VDD#126	XI0/XI1/Q#3	1.24354e-18
C2251	XI1/XI1/D#17	XI1/XI1/XI4/net24#4	3.52091e-17
C2252	XI3/XI1/XI4/PHINOT#9	VDD	4.78049e-18
C2253	XI3/XI1/D#4	PHI#22	1.07136e-17
C2254	SOUT1#20	XI1/XI0/XI1/net2	2.16801e-17
C2255	XI0/XI1/XI4/PHINOT#6	XI0/XI1/XI4/PHINOT#7	4.46757e-18
C2256	XI3/XI1/XI4/PHINOT#4	VDD	2.14306e-17
C2257	XI2/XI1/D#14	RST#8	5.02859e-17
C2258	VDD#160	XI1/XI0/XI0/ANOT	2.05454e-18
C2259	XI0/XI1/D#20	XI0/XI1/D#4	9.89326e-18
C2260	GND#32	GND#31	7.9864e-18
C2261	GND#140	XI1/XI1/D	2.42413e-18
C2262	XI2/XI0/XI0/ANOT#6	net14#3	5.33566e-18
C2263	XI3/XI1/D#10	VDD	1.26139e-17
C2264	XI3/XI1/XI4/net24#11	PHI#23	1.50188e-17
C2265	net7#8	XI1/XI0/XI0/BNOT#14	8.83203e-18
C2266	net7#17	SOUT1#5	2.7909e-17
C2267	XI1/XI1/XI4/net24#11	VDD#123	1.56401e-17
C2268	XI2/XI1/D#17	XI2/XI1/XI4/net24#12	8.08047e-18
C2269	VDD#10	CIN#11	2.54235e-17
C2270	XI2/XI0/XI1/net2#16	SOUT2#5	2.87586e-18
C2271	VDD#130	PHI#4	4.96959e-18
C2272	XI1/XI1/D#19	XI1/XI1/XI4/net24#6	1.52492e-17
C2273	XI1/XI1/Q#11	PHI#12	1.32498e-17
C2274	VDD#78	XI2/XI0/XI0/BNOT#4	1.39714e-18
C2275	SOUT1#14	SOUT1	3.64962e-17
C2276	COUT#5	XI3/XI0/XI1/net2#2	1.85354e-18
C2277	XI1/XI0/XI1/net2#15	net14#10	6.82353e-18
C2278	RST#8	XI2/XI1/D#6	1.04408e-17
C2279	SOUT2#6	net14#5	3.39838e-18
C2280	VDD#155	GND#135	1.78524e-17
C2281	GND#70	PHI#21	5.08165e-18
C2282	XI2/XI0/XI0/BNOT#7	XI2/XI0/XI0/ANOT#9	4.40775e-18
C2283	VDD#70	XI2/XI1/XI4/net24#11	6.32412e-17
C2284	XI2/XI1/D#15	net14#17	5.95074e-18
C2285	XI0/XI1/D	XI0/XI1/XI4/net24#3	2.52567e-18
C2286	XI0/XI1/D#17	PHI#6	1.97458e-18
C2287	XI2/XI1/XI4/net24#11	PHI#16	7.57347e-18
C2288	net21#17	VDD#140	6.83507e-18
C2289	VDD#148	XI2/XI0/XI1/net2#15	3.53013e-18
C2290	XI1/XI1/Q#6	XI1/XI1/D#20	8.17481e-17
C2291	XI2/XI0/XI1/net2#13	RST#8	2.21589e-17
C2292	VDD#142	VDD	1.8633e-17
C2293	net21#14	GND#128	1.08364e-16
C2294	XI0/net1#4	CIN#6	1.35025e-17
C2295	XI0/XI1/Q#9	XI0/XI1/Q#3	2.18451e-18
C2296	XI3/XI0/XI0/ANOT	net21#7	1.29274e-18
C2297	SOUT1#22	net14#21	1.19989e-16
C2298	XI1/XI0/XI1/net2#15	XI1/XI0/XI1/net2#2	6.41939e-18
C2299	SOUT2#18	VDD#112	2.18537e-17
C2300	XI2/net1#4	VDD#76	8.38893e-18
C2301	XI3/XI0/XI0/ANOT#9	net21#3	1.29853e-18
C2302	SOUT2#8	SOUT2#11	8.1418e-18
C2303	VDD#46	XI1/XI0/XI1/net2#3	1.01229e-18
C2304	VDD#86	XI3/XI0/XI0/BNOT#5	5.45774e-17
C2305	XI0/net1#4	XI0/XI0/XI1/net2#3	1.41355e-18
C2306	GND#42	net14#12	4.0234e-17
C2307	XI2/net1#9	XI2/XI0/XI0/BNOT#14	1.07711e-17
C2308	XI1/XI1/Q#6	PHI#11	4.16718e-17
C2309	XI0/XI0/XI1/net2#15	CIN#5	7.43893e-18
C2310	SOUT3#16	SOUT3#19	1.38255e-17
C2311	RST#8	GND#138	7.91186e-18
C2312	XI0/XI0/XI1/net2#15	XI0/XI0/XI1/net2#2	6.41939e-18
C2313	SOUT1#20	XI1/XI0/XI1/net2#3	1.51276e-18
C2314	GND#152	XI0/XI1/XI4/PHINOT#6	1.36671e-17
C2315	XI3/XI0/XI1/net2#13	COUT#3	3.2914e-18
C2316	XI2/XI0/XI0/BNOT#2	XI2/XI0/XI0/BNOT#9	1.3821e-17
C2317	GND#100	XI2/net1#16	9.27251e-18
C2318	GND#28	XI1/XI0/XI0/ANOT#9	5.65589e-18
C2319	VDD#159	SOUT1#20	2.94846e-18
C2320	VDD#22	XI0/XI1/Q	4.68876e-18
C2321	RST#13	XI3/XI0/XI1/net2	1.47319e-17
C2322	XI3/XI0/XI0/BNOT#5	VDD	8.81368e-18
C2323	SOUT3#5	RST#11	3.72778e-17
C2324	XI2/XI1/D#2	XI2/XI1/XI4/net24#2	4.04498e-17
C2325	GND#115	XI0/XI0/XI0/ANOT#3	4.34667e-18
C2326	SOUT0#22	XI0/XI0/XI0/BNOT#4	3.05405e-18
C2327	VDD#2	VDD	1.49508e-17
C2328	VDD#102	SOUT3#20	4.21807e-18
C2329	VDD#141	VDD	1.94359e-17
C2330	XI1/net1#2	SOUT1#6	1.96305e-17
C2331	GND#58	XI2/XI0/XI0/ANOT#3	2.55369e-18
C2332	SOUT0#16	SOUT0#19	1.38255e-17
C2333	SOUT1	VDD#119	1.57577e-17
C2334	GND#101	XI2/XI0/XI0/BNOT#2	3.63595e-18
C2335	VDD#176	VDD	1.01216e-16
C2336	GND#109	SOUT1#3	5.38904e-18
C2337	XI2/XI1/D#17	XI2/XI1/XI4/PHINOT#3	8.962e-19
C2338	XI3/XI1/Q#12	XI3/XI1/XI4/PHINOT#2	2.90831e-18
C2339	VDD#40	VDD#44	3.93119e-17
C2340	XI1/XI0/XI1/net2#13	GND#42	1.11306e-17
C2341	XI3/XI1/D#20	XI3/XI1/XI4/net24#12	1.97297e-17
C2342	VDD#155	XI1/XI0/XI1/net2#2	1.25381e-18
C2343	XI0/XI1/Q#6	VDD#130	1.9494e-18
C2344	GND#123	XI3/XI1/XI4/net24#6	1.96676e-17
C2345	XI3/XI1/D#3	PHI#22	5.34502e-17
C2346	XI1/XI0/XI1/net2#16	XI1/XI0/XI1/net2#15	7.06182e-18
C2347	XI0/XI1/D#15	CIN#11	5.95074e-18
C2348	net21#19	VDD	7.38122e-18
C2349	XI0/XI0/XI0/ANOT#6	GND#6	1.48844e-17
C2350	VDD#24	SOUT0#20	4.21807e-18
C2351	SOUT1#11	XI1/XI0/XI0/ANOT#2	1.22267e-18
C2352	XI2/XI1/Q#6	PHI#17	4.16718e-17
C2353	GND#8	XI0/net1	4.05515e-18
C2354	XI2/XI1/XI4/PHINOT#3	XI2/XI1/D	3.80638e-17
C2355	XI0/XI1/D#10	XI0/net1#2	7.8648e-18
C2356	RST#11	GND#64	1.13456e-17
C2357	SOUT3#11	XI3/XI0/XI0/ANOT#2	1.22267e-18
C2358	net21#17	VDD	6.33291e-18
C2359	GND#132	XI2/XI1/D#2	3.24657e-18
C2360	XI2/XI1/Q#9	SOUT2#16	1.50594e-18
C2361	SOUT0#20	RST#2	1.76518e-17
C2362	CIN#2	VDD#2	3.99391e-18
C2363	VDD#4	VDD	1.68456e-17
C2364	XI3/net1#16	XI3/XI0/XI0/BNOT#9	1.54391e-17
C2365	XI1/net1#9	VDD#52	2.27772e-18
C2366	XI3/net1#9	VDD#138	3.67621e-17
C2367	XI2/XI0/XI0/ANOT#9	net14#3	1.29853e-18
C2368	SOUT2#7	XI2/XI0/XI0/ANOT	5.39732e-17
C2369	XI0/XI1/Q#7	XI0/XI1/XI4/PHINOT	1.21362e-17
C2370	GND#128	RST#11	2.41904e-17
C2371	RST#8	net14#12	7.49192e-18
C2372	PHI#17	VDD#74	5.40385e-18
C2373	VDD#62	XI2/net1#2	1.39754e-17
C2374	XI1/XI0/XI1/net2#16	SOUT1#6	5.16806e-18
C2375	VDD#132	VDD	1.05544e-16
C2376	GND#34	XI1/XI1/D	3.7665e-18
C2377	net21	SOUT3#2	2.69766e-18
C2378	VDD#92	XI3/XI1/XI4/net24#13	1.09794e-18
C2379	SOUT3#24	XI3/XI0/XI0/ANOT#3	2.93467e-18
C2380	XI0/XI1/D#6	RST#1	5.54809e-18
C2381	VDD#40	XI1/XI1/XI4/net24	6.41722e-18
C2382	VDD#5	VDD	2.11985e-17
C2383	SOUT1#7	XI1/XI0/XI0/ANOT	5.39732e-17
C2384	SOUT2#16	SOUT2#17	4.09771e-18
C2385	VDD#140	VDD	2.56909e-17
C2386	RST#8	GND#130	6.19589e-18
C2387	SOUT3	VDD	1.56965e-17
C2388	XI1/XI1/D#19	GND#34	2.48425e-18
C2389	VDD#68	XI2/XI0/XI0/ANOT	4.13602e-18
C2390	XI1/XI1/Q#9	XI1/XI1/Q#8	3.3441e-18
C2391	XI2/XI1/D#17	XI2/XI1/XI4/net24#4	3.52091e-17
C2392	SOUT0#10	XI0/XI0/XI0/BNOT#4	2.61929e-18
C2393	GND#74	GND#73	7.83801e-18
C2394	SOUT2	VDD	1.56965e-17
C2395	VDD#42	XI1/net1#9	2.69821e-18
C2396	GND#147	XI0/XI0/XI1/net2	2.76367e-18
C2397	VDD#162	XI1/net1#2	9.35443e-18
C2398	VDD#119	XI1/XI1/Q#3	1.24354e-18
C2399	XI3/XI1/Q#11	XI3/XI1/Q#2	3.35663e-18
C2400	SOUT1	VDD	1.56965e-17
C2401	XI1/XI0/XI1/net2#13	net7#4	2.31785e-18
C2402	SOUT2#14	SOUT2#15	6.95608e-18
C2403	XI0/XI0/XI0/ANOT#4	VDD	9.31981e-18
C2404	RST#2	GND#10	1.18488e-17
C2405	VDD#129	XI0/XI1/Q	4.97335e-18
C2406	XI1/XI1/XI4/net24#13	XI1/XI1/XI4/net24#2	1.71266e-17
C2407	GND#44	GND#43	7.74457e-18
C2408	SOUT0	VDD	1.56965e-17
C2409	XI1/XI1/XI4/net24#12	SOUT1#19	5.54297e-18
C2410	XI3/XI0/XI0/ANOT#4	XI3/XI0/XI0/BNOT#5	1.1098e-17
C2411	XI3/XI0/XI0/BNOT#9	XI3/XI0/XI0/ANOT#2	4.19591e-17
C2412	XI1/XI0/XI0/BNOT#4	net7#7	2.43471e-17
C2413	SOUT2#10	XI2/XI0/XI0/BNOT#11	3.84272e-17
C2414	XI2/XI1/D#19	XI2/XI1/XI4/net24#6	1.52492e-17
C2415	SOUT2#22	net14#8	5.05993e-18
C2416	GND#107	SOUT1#10	7.13064e-18
C2417	VDD#28	XI1/XI0/XI0/ANOT#4	5.51165e-17
C2418	VDD#126	PHI#8	2.63987e-17
C2419	PHI	VDD	2.24988e-17
C2420	XI2/XI0/XI0/BNOT#4	VDD#147	2.37247e-18
C2421	net21#9	SOUT3#9	3.7545e-17
C2422	XI3/XI1/Q#9	SOUT3#19	5.37314e-18
C2423	XI0/XI1/XI4/net24#11	XI0/XI1/D#4	3.45102e-18
C2424	GND#107	GND#44	9.65661e-18
C2425	XI0/XI1/XI4/net24#4	PHI#6	3.61375e-17
C2426	XI0/XI0/XI0/BNOT#9	XI0/XI0/XI0/ANOT#2	4.19591e-17
C2427	SOUT2#14	VDD#115	1.16528e-17
C2428	XI3/XI0/XI0/BNOT#10	SOUT3#2	7.16694e-18
C2429	XI1/XI1/D#14	SOUT1#5	7.88532e-18
C2430	GND#68	XI3/XI0/XI0/ANOT#6	4.05316e-17
C2431	XI3/XI0/XI0/BNOT#5	net21#19	4.10074e-17
C2432	XI0/XI1/XI4/PHINOT#9	VDD	4.78049e-18
C2433	SOUT2#24	XI2/XI0/XI0/ANOT#2	7.14175e-18
C2434	XI2/XI1/XI4/net24#6	XI2/XI1/D#17	1.49998e-18
C2435	XI2/XI1/D#10	RST#9	3.88703e-18
C2436	VDD#18	VDD#130	1.16687e-17
C2437	XI3/XI1/Q#7	VDD	1.11747e-17
C2438	XI2/XI0/XI1/net2#13	XI2/XI0/XI1/net2	2.66668e-18
C2439	net21#3	SOUT3#3	7.17245e-18
C2440	net14#12	net14#13	4.31453e-18
C2441	XI0/net1	SOUT0#5	4.53739e-18
C2442	GND#94	XI3/XI0/XI0/BNOT#2	3.63595e-18
C2443	XI1/XI0/XI0/ANOT#6	net7#3	5.33566e-18
C2444	XI0/XI1/XI4/PHINOT#4	VDD	2.14306e-17
C2445	XI2/XI0/XI0/ANOT#4	VDD#154	1.1119e-17
C2446	XI3/XI1/Q#5	VDD	1.57977e-17
C2447	RST#8	GND#134	1.95518e-17
C2448	XI2/XI1/XI4/net24	XI2/XI1/D#3	2.28624e-18
C2449	XI0/XI1/D#10	VDD	1.26139e-17
C2450	VDD#137	XI3/XI0/XI1/net2#2	4.26212e-18
C2451	PHI#17	XI2/XI1/Q#2	2.73644e-17
C2452	GND#48	PHI#15	5.08165e-18
C2453	GND#125	XI3/XI1/XI4/PHINOT#6	1.36671e-17
C2454	VDD#48	SOUT1#14	5.47763e-17
C2455	XI3/XI1/D#10	RST#12	3.88703e-18
C2456	RST#4	XI1/net1	3.14306e-18
C2457	VDD#138	XI3/XI0/XI0/ANOT	2.05454e-18
C2458	GND#60	XI2/XI1/D#17	1.61841e-17
C2459	SOUT3#14	SOUT3#15	6.95608e-18
C2460	XI0/XI1/XI4/net24#11	XI0/XI1/D#3	3.27281e-18
C2461	SOUT2#20	XI2/XI0/XI1/net2	2.16801e-17
C2462	net21#12	GND#129	1.3363e-17
C2463	net7#21	VDD#167	7.44569e-18
C2464	XI3/XI1/D#20	XI3/XI1/D#4	9.89326e-18
C2465	XI1/XI1/XI5/net13#5	XI1/XI1/XI5/net13#3	1.65252e-17
C2466	XI2/XI0/XI1/net2#5	SOUT2#6	1.13988e-18
C2467	RST#8	XI2/XI0/XI1/net2#12	1.33951e-17
C2468	XI0/XI1/XI5/net13#5	GND#152	1.65357e-17
C2469	GND#124	GND	4.94454e-17
C2470	VDD#175	XI0/XI1/D#7	2.19078e-17
C2471	XI0/net1#11	SOUT0#7	4.09829e-18
C2472	XI3/XI0/XI1/net2#5	VDD	4.80889e-18
C2473	XI1/XI0/XI1/XI0/net13#2	GND#140	6.62433e-18
C2474	XI0/net1#14	SOUT0#9	2.33071e-18
C2475	XI3/XI1/D#12	RST#12	3.8218e-18
C2476	XI0/XI0/XI1/net2#9	XI0/XI0/XI1/net2#5	1.75967e-17
C2477	GND#139	GND	2.93477e-17
C2478	XI3/net1#6	VDD#137	2.08719e-17
C2479	VDD#64	XI2/XI0/XI1/net2#9	5.41649e-17
C2480	GND#101	XI2/net1#18	1.88957e-17
C2481	XI1/XI1/XI5/net13#5	GND#142	2.13809e-18
C2482	XI1/net1#9	XI1/net1#6	2.47068e-17
C2483	XI2/XI1/XI5/net13#5	GND#133	2.13809e-18
C2484	XI0/XI1/XI5/net13#3	XI0/XI1/XI5/net13	1.34019e-18
C2485	XI1/XI1/XI5/net13#5	GND#143	1.65357e-17
C2486	XI3/net1#14	SOUT3#9	2.33071e-18
C2487	XI2/XI0/XI1/XI0/net13#4	GND#131	1.71714e-17
C2488	XI1/XI0/XI1/XI0/net13#4	GND#140	1.71714e-17
C2489	XI1/net1#6	VDD	9.42787e-18
C2490	XI2/XI1/D#12	RST#9	3.8218e-18
C2491	XI2/net1#11	XI2/net1#9	3.22415e-17
C2492	XI1/XI0/XI1/net2#5	net7#6	4.5401e-18
C2493	SOUT0#11	XI0/net1#11	2.71623e-17
C2494	XI0/XI1/XI5/net13#5	GND#151	2.13809e-18
C2495	XI1/XI1/XI5/net13#3	RST#4	9.65375e-19
C2496	XI3/XI0/XI0/BNOT#14	XI3/net1#6	2.48409e-17
C2497	XI2/XI0/XI1/XI0/net13#4	XI2/XI0/XI1/XI0/net13#2
+ 1.65252e-17
C2498	XI3/XI1/XI5/net13#5	GND#124	2.13809e-18
C2499	GND#72	GND	8.45704e-18
C2500	XI1/XI1/XI5/net13#3	GND#142	1.99937e-17
C2501	GND#95	GND	7.7752e-17
C2502	XI3/XI1/XI5/net13#5	XI3/XI1/D#16	5.59845e-19
C2503	XI2/net1#6	VDD#148	2.08719e-17
C2504	XI2/net1#16	XI2/net1#14	1.21577e-17
C2505	XI0/XI0/XI1/XI0/net13#4	XI0/XI0/XI1/XI0/net13#5
+ 1.39985e-18
C2506	XI1/XI0/XI1/net2#12	SOUT1#5	1.10754e-18
C2507	RST#5	XI1/XI0/XI1/net2#12	1.33951e-17
C2508	XI1/XI1/D#7	XI1/net1#3	3.56068e-18
C2509	XI2/XI1/XI5/net13#5	GND#134	1.65357e-17
C2510	XI1/XI0/XI1/XI0/net13#4	XI1/XI0/XI1/XI0/net13#5
+ 1.39985e-18
C2511	RST#5	XI1/XI0/XI1/XI0/net13#2	1.6172e-17
C2512	VDD#160	XI1/XI0/XI1/net2#5	7.24405e-18
C2513	XI3/net1#18	XI3/XI0/XI0/ANOT#3	4.06446e-18
C2514	XI3/XI0/XI1/net2#12	GND#86	4.27393e-18
C2515	GND#36	GND	1.6487e-17
C2516	XI1/XI1/D#12	VDD	1.03077e-17
C2517	XI3/net1#6	XI3/XI0/XI0/BNOT#3	4.16658e-18
C2518	GND#32	XI1/XI0/XI1/XI0/net13#4	5.09649e-17
C2519	XI0/XI0/XI1/net2#12	GND#148	2.09632e-17
C2520	GND#108	GND	1.00957e-16
C2521	XI2/XI1/D#12	XI2/XI1/D#10	3.30206e-17
C2522	RST#2	XI0/XI0/XI1/XI0/net13#2	1.6172e-17
C2523	XI2/XI0/XI1/net2#9	XI2/XI0/XI1/net2#5	1.75967e-17
C2524	GND#107	XI1/net1#14	2.13647e-17
C2525	XI0/net1#11	XI0/net1#10	1.44781e-17
C2526	XI2/XI0/XI1/net2#9	SOUT2#6	3.59424e-18
C2527	GND#140	GND	1.33841e-17
C2528	XI0/XI1/D#12	RST#3	3.8218e-18
C2529	RST#2	XI0/XI1/XI5/net13#5	1.58559e-17
C2530	XI2/net1#6	XI2/net1#7	1.46041e-17
C2531	XI3/XI0/XI1/XI0/net13#2	RST#11	1.6172e-17
C2532	XI3/net1#18	GND#94	1.88957e-17
C2533	XI1/net1#14	net7#9	4.12965e-18
C2534	GND#70	GND	2.90341e-17
C2535	XI2/XI0/XI1/net2#12	XI2/XI0/XI1/net2#13	2.34768e-17
C2536	XI3/net1#18	XI3/net1#17	4.03534e-18
C2537	GND#126	GND	5.69811e-17
C2538	VDD#161	XI1/XI0/XI1/net2#5	1.30927e-17
C2539	GND#125	GND	6.11034e-17
C2540	XI2/XI0/XI0/BNOT#14	XI2/net1#6	2.48409e-17
C2541	GND#97	GND	7.0778e-17
C2542	XI1/XI0/XI1/net2#5	VDD	4.80889e-18
C2543	XI2/XI0/XI1/net2#12	GND#130	2.09632e-17
C2544	XI2/net1#6	VDD#78	6.13643e-17
C2545	XI2/net1#6	XI2/XI0/XI0/BNOT#3	4.16658e-18
C2546	GND#141	GND	2.21981e-17
C2547	XI1/XI0/XI1/net2#12	GND#42	4.27393e-18
C2548	XI3/XI1/XI5/net13#5	GND#125	1.65357e-17
C2549	GND#68	GND	2.72738e-17
C2550	XI1/XI0/XI1/net2#12	XI1/XI0/XI1/net2#13	2.34768e-17
C2551	XI3/XI0/XI1/net2#5	XI3/net1#4	2.59338e-17
C2552	RST#5	XI1/XI1/XI5/net13#3	1.58114e-17
C2553	GND#96	GND	8.68581e-17
C2554	XI3/net1#11	VDD#138	1.92499e-17
C2555	XI3/XI0/XI1/net2#12	RST#11	1.33951e-17
C2556	GND#128	GND	6.1091e-17
C2557	XI0/XI0/XI1/net2#5	VDD#20	5.77198e-17
C2558	XI1/XI1/XI5/net13#3	XI1/XI1/XI5/net13	1.34019e-18
C2559	XI3/net1#11	XI3/net1#10	1.44781e-17
C2560	XI3/net1#11	VDD	7.88116e-18
C2561	GND#99	GND	9.60155e-17
C2562	XI2/net1#18	XI2/XI0/XI0/ANOT#3	4.06446e-18
C2563	XI2/net1#11	XI2/XI0/XI0/ANOT	7.57752e-18
C2564	GND#142	GND	4.94454e-17
C2565	XI1/XI1/D#12	XI1/XI1/D#11	2.72982e-18
C2566	XI2/XI0/XI1/net2#9	VDD#150	1.45156e-17
C2567	VDD#31	XI1/XI1/D#12	5.07499e-17
C2568	XI2/XI1/D#12	XI2/XI1/D#7	7.32289e-18
C2569	XI2/net1#14	net14#9	4.12965e-18
C2570	XI0/net1#18	SOUT0#24	2.45041e-17
C2571	XI3/XI1/D#7	XI3/XI1/D#12	7.32289e-18
C2572	XI0/net1#14	GND#22	3.1339e-17
C2573	XI2/net1#14	GND#66	3.1339e-17
C2574	XI2/XI1/XI5/net13#3	GND#133	1.99937e-17
C2575	VDD#94	XI3/net1#11	6.16444e-17
C2576	XI3/XI1/XI5/net13#3	XI3/XI1/XI5/net13	1.34019e-18
C2577	XI2/XI0/XI1/net2#9	net14#5	1.21173e-18
C2578	XI1/net1#6	XI1/net1#7	1.46041e-17
C2579	XI0/net1#14	XI0/net1#13	4.02418e-18
C2580	XI2/XI0/XI1/XI0/net13#2	XI2/XI0/XI1/net2#12	4.69772e-17
C2581	XI1/XI1/XI5/net13#5	RST#5	1.58559e-17
C2582	XI1/XI1/D#12	XI1/XI1/D#7	7.32289e-18
C2583	GND#93	XI3/net1#14	2.13647e-17
C2584	XI2/XI1/XI5/net13#3	RST#7	9.65375e-19
C2585	XI3/XI1/XI5/net13#5	RST#10	3.93763e-18
C2586	XI2/XI0/XI1/net2#5	VDD#72	5.77198e-17
C2587	VDD#140	XI3/XI0/XI1/net2#9	6.37152e-18
C2588	GND#28	GND	8.45704e-18
C2589	XI0/XI1/XI5/net13#3	GND#8	5.09163e-17
C2590	GND#109	GND	7.7752e-17
C2591	XI0/net1#11	VDD#171	1.92499e-17
C2592	XI3/XI1/D#12	XI3/XI1/D#11	2.72982e-18
C2593	XI0/XI1/D#7	VDD#10	5.39472e-17
C2594	GND#66	GND	8.80845e-18
C2595	XI0/XI1/XI5/net13#5	RST#1	3.93763e-18
C2596	XI0/XI0/XI1/net2#9	VDD	5.99038e-18
C2597	XI3/XI0/XI1/net2#12	GND#121	2.09632e-17
C2598	GND#100	GND	7.75707e-17
C2599	XI2/XI1/D#7	VDD	1.03467e-17
C2600	VDD#138	XI3/XI0/XI1/net2#5	7.24405e-18
C2601	net21#8	XI3/net1#6	3.2757e-18
C2602	XI3/XI1/D#7	XI3/XI1/D#8	2.66591e-18
C2603	XI0/XI1/D#12	XI0/XI1/D#7	7.32289e-18
C2604	XI3/XI0/XI1/XI0/net13#2	GND#122	6.62433e-18
C2605	XI0/XI1/XI5/net13#3	GND#151	1.99937e-17
C2606	XI0/XI0/XI1/net2#9	SOUT0#6	3.59424e-18
C2607	XI1/XI0/XI1/net2#12	net7#4	3.76602e-18
C2608	XI0/net1#6	CIN#7	7.64271e-18
C2609	XI2/net1#14	XI2/net1#13	4.02418e-18
C2610	XI3/XI1/XI5/net13#3	GND#74	5.09163e-17
C2611	XI2/XI1/XI5/net13#5	XI2/XI1/XI5/net13#3	1.65252e-17
C2612	XI1/net1#6	XI1/XI0/XI0/BNOT#3	4.16658e-18
C2613	XI3/net1#14	SOUT3#10	1.90893e-17
C2614	GND#135	GND	5.69811e-17
C2615	GND#129	GND	4.55207e-17
C2616	XI3/XI1/D#7	VDD#88	5.39472e-17
C2617	GND#104	GND	7.0778e-17
C2618	XI3/net1#16	XI3/net1#14	1.21577e-17
C2619	CIN#8	XI0/net1#11	2.44833e-18
C2620	XI2/XI0/XI1/net2#9	XI2/net1#4	1.93606e-17
C2621	XI2/XI0/XI1/net2#12	XI2/XI0/XI1/net2	9.43555e-19
C2622	VDD#16	XI0/net1#11	6.16444e-17
C2623	VDD#161	XI1/XI0/XI1/net2#9	1.45156e-17
C2624	XI2/net1#6	net14#7	7.64271e-18
C2625	net7#8	XI1/net1#11	2.44833e-18
C2626	XI0/XI1/D#7	XI0/net1#3	3.56068e-18
C2627	XI0/net1#18	XI0/net1#17	4.03534e-18
C2628	XI3/XI0/XI1/net2#9	net21#5	1.21173e-18
C2629	XI0/XI1/D#6	XI0/XI1/XI5/net13#5	5.14071e-17
C2630	XI1/net1#11	VDD	7.88116e-18
C2631	XI3/XI0/XI1/net2#9	VDD	5.99038e-18
C2632	GND#26	GND	2.90341e-17
C2633	GND#143	GND	6.11034e-17
C2634	XI3/XI0/XI1/net2#9	XI3/net1#4	1.93606e-17
C2635	XI1/net1#14	SOUT1#9	2.33071e-18
C2636	XI2/net1#18	SOUT2#24	2.45041e-17
C2637	XI0/net1#6	VDD#170	2.08719e-17
C2638	VDD#150	XI2/XI0/XI1/net2#5	1.30927e-17
C2639	XI2/net1#14	SOUT2#9	2.33071e-18
C2640	XI2/XI1/D#15	XI2/XI1/XI5/net13#5	1.42469e-18
C2641	XI1/net1#18	XI1/net1#14	2.75871e-18
C2642	XI2/XI0/XI1/net2#5	XI2/XI0/XI1/net2#4	1.50642e-18
C2643	XI3/net1#18	XI3/XI0/XI0/BNOT#2	2.19446e-18
C2644	XI2/net1#18	XI2/net1#14	2.75871e-18
C2645	XI0/XI0/XI1/net2#12	XI0/XI0/XI1/net2	9.43555e-19
C2646	XI0/XI1/XI5/net13#5	XI0/XI1/D#15	1.42469e-18
C2647	XI3/XI0/XI1/XI0/net13#4	RST#11	1.62165e-17
C2648	GND#24	GND	2.72738e-17
C2649	GND#110	GND	8.68581e-17
C2650	XI1/net1#18	XI1/XI0/XI0/BNOT	2.2742e-18
C2651	XI3/XI0/XI1/net2#12	SOUT3#5	1.10754e-18
C2652	XI3/XI1/D#12	XI3/XI1/D#10	3.30206e-17
C2653	XI1/XI0/XI1/XI0/net13#4	XI1/XI0/XI1/XI0/net13#2
+ 1.65252e-17
C2654	GND#146	GND	6.1091e-17
C2655	GND#113	GND	9.60155e-17
C2656	XI2/net1#6	VDD	9.42787e-18
C2657	XI3/net1#11	XI3/net1#9	3.22415e-17
C2658	XI1/XI1/D#6	XI1/XI1/XI5/net13#5	5.14071e-17
C2659	XI2/net1#18	XI2/XI0/XI0/BNOT#2	2.19446e-18
C2660	XI0/XI0/XI1/XI0/net13#2	GND#149	6.62433e-18
C2661	XI1/XI1/XI5/net13#5	XI1/XI1/XI5/net13#4	1.49662e-18
C2662	XI1/XI0/XI1/net2#9	net7#5	1.21173e-18
C2663	XI0/net1#11	XI0/net1#9	3.22415e-17
C2664	GND#130	GND	2.93477e-17
C2665	XI3/XI0/XI1/XI0/net13#4	GND#122	1.71714e-17
C2666	XI0/XI1/D#12	XI0/XI1/D#11	2.72982e-18
C2667	XI1/XI0/XI1/net2#12	GND#139	2.09632e-17
C2668	XI2/XI0/XI1/XI0/net13#2	RST#8	1.6172e-17
C2669	XI0/net1#18	XI0/XI0/XI0/ANOT#3	4.06446e-18
C2670	XI3/XI0/XI1/net2#5	net21#6	4.5401e-18
C2671	XI0/XI0/XI1/XI0/net13#4	GND#149	1.71714e-17
C2672	net21#8	XI3/net1#11	2.44833e-18
C2673	VDD#83	XI3/XI1/D#12	5.07499e-17
C2674	RST#2	XI0/XI0/XI1/net2#12	1.33951e-17
C2675	XI0/XI0/XI1/net2#9	XI0/net1#4	1.93606e-17
C2676	XI1/XI0/XI1/net2#9	VDD#162	6.37152e-18
C2677	XI3/XI0/XI1/net2#5	XI3/XI0/XI1/net2#4	1.50642e-18
C2678	net14#8	XI2/net1#6	3.2757e-18
C2679	GND#22	GND	8.80845e-18
C2680	GND#114	GND	7.75707e-17
C2681	XI3/XI1/D#10	XI3/XI1/D#7	3.40394e-17
C2682	GND#144	GND	5.69811e-17
C2683	XI0/XI0/XI1/net2#5	XI0/net1#4	2.59338e-17
C2684	XI3/net1#11	XI3/XI0/XI0/ANOT	7.57752e-18
C2685	GND#111	GND	7.0778e-17
C2686	XI2/XI1/D#12	XI2/XI1/D#11	2.72982e-18
C2687	XI3/XI1/XI5/net13#3	XI3/XI1/D#15	1.98365e-18
C2688	XI1/net1#14	SOUT1#10	1.90893e-17
C2689	GND#58	GND	1.6487e-17
C2690	XI2/XI1/D#6	XI2/XI1/XI5/net13#5	5.14071e-17
C2691	GND#101	GND	1.00957e-16
C2692	XI3/XI0/XI1/net2#9	VDD#139	1.45156e-17
C2693	XI3/XI0/XI1/net2#12	XI3/XI0/XI1/net2#13	2.34768e-17
C2694	GND#147	GND	4.55207e-17
C2695	XI1/net1#6	VDD#159	2.08719e-17
C2696	XI2/XI0/XI1/net2#9	XI2/XI0/XI1/net2#7	1.56189e-18
C2697	XI2/net1#11	VDD#149	1.92499e-17
C2698	XI1/net1#14	XI1/net1#13	4.02418e-18
C2699	XI0/XI0/XI0/BNOT#14	XI0/net1#6	2.48409e-17
C2700	XI2/XI0/XI1/net2#12	XI2/XI0/XI1/net2#10	3.45593e-18
C2701	GND#131	GND	1.33841e-17
C2702	XI2/XI1/D#12	VDD	1.03077e-17
C2703	XI3/XI1/XI5/net13#3	RST#10	9.65375e-19
C2704	GND#14	XI0/net1#18	3.12263e-17
C2705	VDD#171	XI0/XI0/XI1/net2#5	7.24405e-18
C2706	XI0/XI1/D#7	XI0/XI1/D#8	2.66591e-18
C2707	XI0/net1#6	XI0/XI0/XI0/BNOT#3	4.16658e-18
C2708	GND#36	XI1/net1#18	3.12263e-17
C2709	VDD#153	XI2/XI1/D#7	2.19078e-17
C2710	XI1/XI0/XI1/net2#9	XI1/XI0/XI1/net2#5	1.75967e-17
C2711	SOUT3#11	XI3/net1#11	2.71623e-17
C2712	XI1/net1#6	XI1/net1#11	4.94255e-18
C2713	XI0/XI1/XI5/net13#5	XI0/XI1/XI5/net13#4	1.49662e-18
C2714	XI0/net1#18	XI0/net1#16	1.59717e-17
C2715	RST#11	XI3/XI1/XI5/net13#5	1.58559e-17
C2716	XI0/XI0/XI1/net2#5	SOUT0#6	1.13988e-18
C2717	XI2/XI0/XI1/XI0/net13#2	XI2/XI0/XI1/XI0/net13	1.47724e-18
C2718	GND#132	GND	2.21981e-17
C2719	XI0/net1#11	XI0/net1#6	4.94255e-18
C2720	XI3/net1#18	XI3/XI0/XI0/BNOT	2.2742e-18
C2721	XI2/net1#6	XI2/net1#11	4.94255e-18
C2722	XI0/XI1/D#7	VDD	1.03467e-17
C2723	VDD#164	XI1/XI1/D#7	2.19078e-17
C2724	XI2/XI0/XI1/net2#5	VDD	4.80889e-18
C2725	XI1/XI0/XI1/XI0/net13#2	XI1/XI0/XI1/net2#12	4.69772e-17
C2726	XI0/net1#18	XI0/XI0/XI0/BNOT#2	2.19446e-18
C2727	GND#114	XI0/net1#14	2.13647e-17
C2728	XI3/net1#6	XI3/net1#7	1.46041e-17
C2729	VDD#139	XI3/XI0/XI1/net2#5	1.30927e-17
C2730	XI2/XI1/XI5/net13#5	RST#7	3.93763e-18
C2731	XI1/net1#11	XI1/XI0/XI0/ANOT	7.57752e-18
C2732	GND#58	XI2/net1#18	3.12263e-17
C2733	XI2/XI0/XI1/net2#12	SOUT2#5	1.10754e-18
C2734	XI3/net1#14	XI3/net1#13	4.02418e-18
C2735	XI1/XI1/XI5/net13#5	RST#4	3.93763e-18
C2736	GND#119	GND	6.10818e-17
C2737	VDD#42	XI1/net1#11	6.16444e-17
C2738	XI1/net1#18	XI1/net1#16	1.59717e-17
C2739	XI0/XI0/XI1/net2#12	XI0/XI0/XI1/net2#13	2.34768e-17
C2740	GND#92	GND	9.61308e-17
C2741	GND#133	GND	4.94454e-17
C2742	VDD#143	XI3/XI1/D#12	1.34081e-17
C2743	XI3/XI1/XI5/net13#3	RST#11	1.58114e-17
C2744	XI3/net1#11	XI3/net1#6	4.94255e-18
C2745	GND#148	GND	2.93477e-17
C2746	XI3/XI1/D#6	XI3/XI1/XI5/net13#5	5.14071e-17
C2747	XI0/net1#14	SOUT0#10	1.90893e-17
C2748	XI1/XI0/XI1/net2#9	VDD	5.99038e-18
C2749	XI3/XI1/XI5/net13#5	XI3/XI1/XI5/net13#4	1.49662e-18
C2750	XI2/net1#11	SOUT2#7	4.09829e-18
C2751	XI0/XI1/D#12	XI0/XI1/D#10	3.30206e-17
C2752	XI1/XI0/XI0/BNOT#14	XI1/net1#6	2.48409e-17
C2753	XI2/net1#18	XI2/XI0/XI0/BNOT	2.2742e-18
C2754	XI3/XI0/XI1/net2#12	net21#4	3.76602e-18
C2755	XI1/net1#11	XI1/net1#10	1.44781e-17
C2756	XI3/XI1/D#7	VDD	1.03467e-17
C2757	XI2/XI0/XI1/XI0/net13#2	GND#131	6.62433e-18
C2758	XI2/net1#9	XI2/net1#6	2.47068e-17
C2759	XI1/XI1/D#10	XI1/XI1/D#7	3.40394e-17
C2760	XI0/XI0/XI1/net2#5	XI0/XI0/XI1/net2#4	1.50642e-18
C2761	VDD#5	XI0/XI1/D#12	5.07499e-17
C2762	XI3/XI1/XI5/net13#5	XI3/XI1/XI5/net13#3	1.65252e-17
C2763	XI1/XI1/XI5/net13#3	XI1/XI1/D#15	1.98365e-18
C2764	XI3/XI0/XI1/net2#9	SOUT3#6	3.59424e-18
C2765	XI3/XI0/XI1/XI0/net13#2	GND#121	1.2558e-17
C2766	XI3/net1#9	XI3/net1#6	2.47068e-17
C2767	XI0/net1#11	XI0/XI0/XI0/ANOT	7.57752e-18
C2768	VDD#173	XI0/XI0/XI1/net2#9	6.37152e-18
C2769	XI0/XI0/XI1/net2#12	XI0/XI0/XI1/net2#10	3.45593e-18
C2770	GND#80	XI3/net1#18	3.12263e-17
C2771	GND#50	GND	8.45704e-18
C2772	XI2/XI0/XI1/net2#9	VDD#151	6.37152e-18
C2773	XI0/XI1/D#12	VDD	1.03077e-17
C2774	XI2/net1#11	XI2/net1#10	1.44781e-17
C2775	XI0/net1#16	XI0/net1#14	1.21577e-17
C2776	XI2/net1#14	GND#100	2.13647e-17
C2777	XI1/XI0/XI1/net2#9	SOUT1#6	3.59424e-18
C2778	XI2/net1#18	XI2/net1#16	1.59717e-17
C2779	XI0/XI1/XI5/net13#5	XI0/XI1/D#16	5.59845e-19
C2780	GND#102	GND	7.7752e-17
C2781	CIN#8	XI0/net1#6	3.2757e-18
C2782	GND#88	GND	8.80845e-18
C2783	VDD#149	XI2/XI0/XI1/net2#5	7.24405e-18
C2784	VDD#38	XI1/XI0/XI1/net2#9	5.41649e-17
C2785	XI2/XI0/XI1/XI0/net13#4	XI2/XI0/XI1/XI0/net13#5
+ 1.39985e-18
C2786	GND#93	GND	7.75707e-17
C2787	RST#5	XI1/XI0/XI1/XI0/net13#4	1.62165e-17
C2788	XI1/XI0/XI1/net2#5	XI1/net1#4	2.59338e-17
C2789	XI0/net1#6	VDD	9.42787e-18
C2790	XI1/XI0/XI1/net2#9	XI1/net1#4	1.93606e-17
C2791	XI0/net1#18	XI0/net1#14	2.75871e-18
C2792	SOUT2#11	XI2/net1#11	2.71623e-17
C2793	GND#14	GND	1.6487e-17
C2794	XI3/XI0/XI1/net2#9	XI3/XI0/XI1/net2#5	1.75967e-17
C2795	GND#115	GND	9.19313e-17
C2796	net14#8	XI2/net1#11	2.44833e-18
C2797	XI2/net1#18	XI2/net1#17	4.03534e-18
C2798	XI2/XI1/D#12	VDD#154	1.34081e-17
C2799	XI0/XI1/XI5/net13#3	XI0/XI1/XI5/net13#5	1.65252e-17
C2800	XI0/XI0/XI1/net2#9	XI0/XI0/XI1/net2#7	1.56189e-18
C2801	XI3/net1#18	XI3/net1#14	2.75871e-18
C2802	XI3/XI0/XI1/XI0/net13#2	XI3/XI0/XI1/XI0/net13	1.47724e-18
C2803	XI1/XI0/XI1/net2#5	VDD#46	5.77198e-17
C2804	GND#120	GND	4.55382e-17
C2805	XI1/net1#11	XI1/net1#9	3.22415e-17
C2806	XI1/net1#14	GND#44	3.1339e-17
C2807	GND#149	GND	1.33841e-17
C2808	XI2/net1#14	SOUT2#10	1.90893e-17
C2809	VDD#12	XI0/XI0/XI1/net2#9	5.41649e-17
C2810	XI3/XI0/XI1/net2#5	SOUT3#6	1.13988e-18
C2811	XI2/XI1/XI5/net13#5	RST#8	1.58559e-17
C2812	XI0/XI0/XI1/net2#5	VDD	4.80889e-18
C2813	XI0/net1#14	CIN#9	4.12965e-18
C2814	XI2/XI0/XI1/XI0/net13#2	GND#130	1.2558e-17
C2815	GND#48	GND	2.90341e-17
C2816	GND#54	XI2/XI0/XI1/XI0/net13#4	5.09649e-17
C2817	XI1/XI1/D#12	RST#6	3.8218e-18
C2818	GND#134	GND	6.11034e-17
C2819	XI0/XI0/XI1/XI0/net13#4	XI0/XI0/XI1/XI0/net13#2
+ 1.65252e-17
C2820	XI1/XI0/XI1/net2#5	XI1/XI0/XI1/net2#4	1.50642e-18
C2821	RST#8	XI2/XI1/XI5/net13#3	1.58114e-17
C2822	XI3/net1#6	VDD	9.42787e-18
C2823	XI3/XI0/XI1/XI0/net13#4	XI3/XI0/XI1/XI0/net13#2
+ 1.65252e-17
C2824	GND#150	GND	2.21981e-17
C2825	RST#2	XI0/XI0/XI1/XI0/net13#4	1.62165e-17
C2826	XI3/net1#18	XI3/net1#16	1.59717e-17
C2827	XI0/XI0/XI1/net2#12	CIN#4	3.76602e-18
C2828	XI2/net1#11	VDD	7.88116e-18
C2829	XI1/net1#18	XI1/net1#17	4.03534e-18
C2830	XI2/XI1/XI5/net13#5	XI2/XI1/XI5/net13#4	1.49662e-18
C2831	XI3/XI0/XI1/net2#9	XI3/XI0/XI1/net2#7	1.56189e-18
C2832	XI1/net1#6	net7#7	7.64271e-18
C2833	GND#46	GND	2.72738e-17
C2834	XI1/net1#18	SOUT1#24	2.45041e-17
C2835	XI3/net1#14	GND#88	3.1339e-17
C2836	VDD#90	XI3/XI0/XI1/net2#9	5.41649e-17
C2837	XI1/XI1/XI5/net13#5	XI1/XI1/D#16	5.59845e-19
C2838	GND#103	GND	8.68581e-17
C2839	XI0/XI0/XI1/XI0/net13#2	XI0/XI0/XI1/XI0/net13	1.47724e-18
C2840	XI3/XI1/XI5/net13#3	GND#124	1.99937e-17
C2841	GND#76	XI3/XI0/XI1/XI0/net13#4	5.09649e-17
C2842	GND#137	GND	6.1091e-17
C2843	XI0/net1#18	XI0/XI0/XI0/BNOT	2.2742e-18
C2844	GND#106	GND	9.60155e-17
C2845	XI1/XI0/XI1/net2#12	XI1/XI0/XI1/net2	9.43555e-19
C2846	XI2/XI1/D#7	XI2/XI1/D#8	2.66591e-18
C2847	GND#151	GND	4.94454e-17
C2848	XI0/XI0/XI1/net2#12	GND#20	4.27393e-18
C2849	XI1/XI0/XI1/net2#12	XI1/XI0/XI1/net2#10	3.45593e-18
C2850	XI3/XI0/XI1/net2#12	XI3/XI0/XI1/net2#10	3.45593e-18
C2851	XI0/net1#9	XI0/net1#6	2.47068e-17
C2852	XI1/net1#18	XI1/XI0/XI0/BNOT#2	2.19446e-18
C2853	XI0/XI1/D#10	XI0/XI1/D#7	3.40394e-17
C2854	VDD#57	XI2/XI1/D#12	5.07499e-17
C2855	XI1/XI0/XI1/net2#9	XI1/XI0/XI1/net2#7	1.56189e-18
C2856	GND#121	GND	2.93302e-17
C2857	VDD#172	XI0/XI0/XI1/net2#9	1.45156e-17
C2858	XI0/XI1/XI5/net13#3	XI0/XI1/D#15	1.98365e-18
C2859	XI3/XI0/XI1/net2#5	VDD#98	5.77198e-17
C2860	VDD#165	XI1/XI1/D#12	1.34081e-17
C2861	XI3/XI0/XI1/XI0/net13#4	XI3/XI0/XI1/XI0/net13#5
+ 1.39985e-18
C2862	XI3/XI1/D#7	XI3/net1#3	3.56068e-18
C2863	GND#10	XI0/XI0/XI1/XI0/net13#4	5.09649e-17
C2864	XI1/XI1/D#15	XI1/XI1/XI5/net13#5	1.42469e-18
C2865	XI1/XI0/XI1/XI0/net13#2	GND#139	1.2558e-17
C2866	XI0/XI0/XI1/net2#12	SOUT0#5	1.10754e-18
C2867	XI1/net1#6	VDD#52	6.13643e-17
C2868	SOUT1#11	XI1/net1#11	2.71623e-17
C2869	XI1/net1#16	XI1/net1#14	1.21577e-17
C2870	XI3/net1#6	VDD#104	6.13643e-17
C2871	XI1/XI1/D#12	XI1/XI1/D#10	3.30206e-17
C2872	GND#6	GND	8.45704e-18
C2873	XI0/XI0/XI1/net2#5	CIN#6	4.5401e-18
C2874	XI2/XI1/D#10	XI2/XI1/D#7	3.40394e-17
C2875	GND#116	GND	4.46754e-17
C2876	XI2/XI1/XI5/net13#3	XI2/XI1/D#15	1.98365e-18
C2877	GND#44	GND	8.80845e-18
C2878	XI1/net1#14	XI1/XI0/XI0/BNOT#11	4.26343e-18
C2879	XI0/XI0/XI1/net2#9	CIN#5	1.21173e-18
C2880	GND#107	GND	7.75707e-17
C2881	XI0/XI0/XI0/BNOT#11	XI0/net1#14	4.26343e-18
C2882	XI1/net1#11	VDD#160	1.92499e-17
C2883	XI1/XI1/XI5/net13#3	GND#30	5.09163e-17
C2884	XI0/XI1/XI5/net13#3	RST#2	1.58114e-17
C2885	XI1/XI1/D#7	XI1/XI1/D#8	2.66591e-18
C2886	XI2/XI0/XI1/XI0/net13#4	RST#8	1.62165e-17
C2887	XI0/net1#18	GND#115	1.88957e-17
C2888	XI1/XI1/D#7	VDD#36	5.39472e-17
C2889	XI3/XI1/XI5/net13#5	XI3/XI1/D#15	1.42469e-18
C2890	XI2/XI0/XI0/BNOT#11	XI2/net1#14	4.26343e-18
C2891	XI2/XI1/XI5/net13#3	GND#52	5.09163e-17
C2892	GND#80	GND	1.6487e-17
C2893	VDD#68	XI2/net1#11	6.16444e-17
C2894	GND#94	GND	1.00957e-16
C2895	XI2/XI1/D#7	VDD#62	5.39472e-17
C2896	XI2/XI0/XI1/net2#5	net14#6	4.5401e-18
C2897	XI2/XI1/XI5/net13#5	XI2/XI1/D#16	5.59845e-19
C2898	XI0/net1#11	VDD	7.88116e-18
C2899	VDD#142	XI3/XI1/D#7	2.19078e-17
C2900	GND#138	GND	4.55207e-17
C2901	XI2/XI0/XI1/net2#5	XI2/net1#4	2.59338e-17
C2902	XI0/net1#6	XI0/net1#7	1.46041e-17
C2903	XI2/XI1/D#7	XI2/net1#3	3.56068e-18
C2904	XI1/XI0/XI1/XI0/net13#2	XI1/XI0/XI1/XI0/net13	1.47724e-18
C2905	XI3/XI0/XI1/XI0/net13#2	XI3/XI0/XI1/net2#12	4.69772e-17
C2906	GND#122	GND	1.33841e-17
C2907	XI2/XI0/XI1/net2#12	net14#4	3.76602e-18
C2908	XI2/XI1/XI5/net13#3	XI2/XI1/XI5/net13	1.34019e-18
C2909	XI1/XI1/D#7	VDD	1.03467e-17
C2910	net7#8	XI1/net1#6	3.2757e-18
C2911	XI3/XI0/XI1/net2#12	XI3/XI0/XI1/net2	9.43555e-19
C2912	XI2/XI0/XI1/net2#12	GND#64	4.27393e-18
C2913	GND#4	GND	2.90341e-17
C2914	XI1/XI0/XI1/net2#5	SOUT1#6	1.13988e-18
C2915	XI0/net1#6	VDD#26	6.13643e-17
C2916	GND#152	GND	8.46488e-17
C2917	XI0/XI1/XI5/net13#3	RST#1	9.65375e-19
C2918	XI3/XI0/XI0/BNOT#11	XI3/net1#14	4.26343e-18
C2919	GND#108	XI1/net1#18	1.88957e-17
C2920	XI3/net1#18	SOUT3#24	2.45041e-17
C2921	XI3/XI1/D#12	VDD	1.03077e-17
C2922	XI0/XI0/XI1/XI0/net13#2	XI0/XI0/XI1/net2#12	4.69772e-17
C2923	XI3/net1#11	SOUT3#7	4.09829e-18
C2924	XI3/net1#6	net21#7	7.64271e-18
C2925	VDD#172	XI0/XI0/XI1/net2#5	1.30927e-17
C2926	GND#123	GND	2.21981e-17
C2927	GND#2	GND	2.72738e-17
C2928	GND#117	GND	1.06311e-16
C2929	GND#89	GND	4.72899e-17
C2930	GND#118	GND	6.87042e-17
C2931	XI1/net1#18	XI1/XI0/XI0/ANOT#3	4.06446e-18
C2932	XI3/net1#14	net21#9	4.12965e-18
C2933	XI2/XI0/XI1/net2#9	VDD	5.99038e-18
C2934	XI0/XI0/XI1/XI0/net13#2	GND#148	1.2558e-17
C2935	GND#90	GND	4.58994e-17
C2936	VDD#176	XI0/XI1/D#12	1.34081e-17
C2937	XI1/net1#11	SOUT1#7	4.09829e-18
C2938	GND#14	CIN#13	6.6296e-19
C2939	GND#20	CIN#4	7.67752e-19
C2940	GND#2	CIN#2	8.17588e-19
C2941	GND#113	CIN#8	1.04902e-18
C2942	XI1/XI1/D#20	XI1/XI1/Q	3.0256e-19
C2943	XI1/XI1/D#17	XI1/XI1/Q#3	3.77893e-19
C2944	XI1/XI1/Q#6	XI1/XI1/D#4	4.04483e-19
C2945	XI1/XI1/Q#5	XI1/XI1/D#3	4.90626e-19
C2946	XI1/XI1/D#17	XI1/XI1/Q#2	5.79029e-19
C2947	XI1/XI1/D#4	XI1/XI1/Q	6.8315e-19
C2948	CIN#11	RST#3	1.2685e-18
C2949	SOUT0#24	CIN#9	5.74591e-19
C2950	CIN#13	SOUT0#11	8.62763e-19
C2951	CIN#13	SOUT0#1	9.73491e-19
C2952	GND#60	PHI#18	1.372e-18
C2953	GND#38	PHI#12	1.372e-18
C2954	GND#16	PHI#6	1.372e-18
C2955	GND#125	PHI#21	3.38517e-18
C2956	GND#134	PHI#15	3.38517e-18
C2957	GND#143	PHI#9	3.38517e-18
C2958	GND#152	PHI#3	3.38517e-18
C2959	VDD#12	CIN#6	4.8046e-19
C2960	CIN#5	VDD	5.05446e-19
C2961	VDD#24	CIN#6	8.61141e-19
C2962	CIN#2	VDD#8	1.30482e-18
C2963	CIN#13	VDD#172	1.41225e-18
C2964	GND#122	RST#11	9.48137e-19
C2965	GND#131	RST#8	9.48137e-19
C2966	GND#140	RST#5	9.48137e-19
C2967	GND#152	RST#1	2.53688e-18
C2968	GND#125	RST#10	2.53688e-18
C2969	GND#134	RST#7	2.53688e-18
C2970	GND#143	RST#4	2.53688e-18
C2971	RST#13	GND#121	3.06476e-18
C2972	RST#11	GND#121	3.10681e-18
C2973	XI0/net1#18	CIN#9	3.7252e-19
C2974	XI0/net1#11	CIN#6	3.75673e-19
C2975	XI0/net1#4	CIN#11	4.08444e-19
C2976	XI0/net1#9	CIN#7	7.33206e-19
C2977	XI0/net1#11	CIN#7	7.62892e-19
C2978	XI0/net1#16	CIN#9	9.2752e-19
C2979	GND#113	SOUT0#9	8.94058e-19
C2980	GND#14	SOUT0#3	1.60329e-18
C2981	XI0/XI1/D#14	CIN#4	1.47002e-18
C2982	GND#106	SOUT1#9	8.94058e-19
C2983	GND#36	SOUT1#3	1.60329e-18
C2984	COUT#7	VDD#104	1.06668e-18
C2985	XI0/XI0/XI0/BNOT#5	CIN#1	9.33843e-19
C2986	XI0/XI0/XI0/BNOT#7	CIN#3	1.29331e-18
C2987	CIN#13	XI0/XI0/XI0/ANOT	6.60017e-19
C2988	XI0/XI0/XI0/ANOT	CIN#8	8.2626e-19
C2989	GND#99	SOUT2#9	8.94058e-19
C2990	GND#58	SOUT2#3	1.60329e-18
C2991	GND#92	SOUT3#9	8.94058e-19
C2992	GND#80	SOUT3#3	1.60329e-18
C2993	GND#119	VDD#105	2.63264e-18
C2994	GND#128	VDD#112	2.63264e-18
C2995	GND#137	VDD#119	2.63264e-18
C2996	GND#146	VDD#126	2.63264e-18
C2997	GND#92	VDD#133	3.85922e-18
C2998	GND#99	VDD#144	3.85922e-18
C2999	GND#106	VDD#155	3.85922e-18
C3000	GND#113	VDD#166	3.85922e-18
C3001	GND#119	VDD	6.08627e-18
C3002	GND#128	VDD	6.08627e-18
C3003	GND#137	VDD	6.08627e-18
C3004	GND#146	VDD	6.08627e-18
C3005	XI1/XI1/XI4/net24#4	XI1/XI1/Q#2	6.00447e-19
C3006	GND#42	net7#4	7.67752e-19
C3007	GND#24	net7#2	8.17588e-19
C3008	GND#106	net7#8	1.04902e-18
C3009	GND#146	net7#12	1.33266e-18
C3010	GND#28	net7#3	1.73249e-18
C3011	GND#44	net7#9	2.55369e-18
C3012	XI1/XI0/XI0/BNOT#14	XI1/XI0/XI0/ANOT	6.36598e-19
C3013	XI1/XI0/XI0/BNOT#11	XI1/XI0/XI0/ANOT#2	7.40945e-19
C3014	VDD#92	PHI#23	1.48609e-18
C3015	VDD#66	PHI#17	1.48609e-18
C3016	VDD#40	PHI#11	1.48609e-18
C3017	VDD#14	PHI#5	1.48609e-18
C3018	VDD#18	PHI#4	2.37746e-18
C3019	VDD#96	PHI#22	2.37746e-18
C3020	VDD#70	PHI#16	2.37746e-18
C3021	VDD#44	PHI#10	2.37746e-18
C3022	VDD#111	PHI#19	4.6061e-18
C3023	VDD#118	PHI#13	4.6061e-18
C3024	VDD#125	PHI#7	4.6061e-18
C3025	VDD#132	PHI#1	4.6061e-18
C3026	XI0/XI1/D#15	GND#151	1.19132e-18
C3027	XI0/XI1/D#14	GND#150	1.22638e-18
C3028	GND#12	XI0/XI1/XI4/net24#3	9.20398e-19
C3029	GND#12	XI0/XI1/XI4/net24#2	9.87977e-19
C3030	GND#113	XI0/XI0/XI0/BNOT#3	6.89259e-19
C3031	GND#113	XI0/XI0/XI0/BNOT#4	7.0191e-19
C3032	XI0/XI1/D#19	PHI#2	8.74572e-19
C3033	GND#147	XI0/XI1/Q#2	4.8289e-19
C3034	VDD#166	SOUT0#20	5.92296e-19
C3035	VDD#10	SOUT0#6	6.94836e-19
C3036	SOUT0#11	VDD#171	7.64293e-19
C3037	SOUT0	VDD#127	7.94421e-19
C3038	VDD#16	SOUT0#1	1.21155e-18
C3039	SOUT0#11	VDD	1.24623e-18
C3040	SOUT0#8	VDD	2.30293e-18
C3041	VDD#174	SOUT0#1	2.33481e-18
C3042	XI0/XI1/XI4/net24#2	PHI#6	7.75967e-19
C3043	XI0/XI1/XI4/net24#2	PHI#5	9.535e-19
C3044	VDD#155	SOUT1#20	5.92296e-19
C3045	VDD#36	SOUT1#6	6.94836e-19
C3046	SOUT1#11	VDD#160	7.64293e-19
C3047	SOUT1	VDD#120	7.94421e-19
C3048	VDD#42	SOUT1#1	1.21155e-18
C3049	SOUT1#11	VDD	1.24623e-18
C3050	SOUT1#8	VDD	2.30293e-18
C3051	VDD#163	SOUT1#1	2.33481e-18
C3052	XI0/XI1/D#15	RST#3	1.25112e-18
C3053	SOUT0#2	XI0/net1#3	5.53224e-19
C3054	XI0/net1#2	SOUT0#1	5.64483e-19
C3055	XI0/net1#3	SOUT0#6	9.94394e-19
C3056	SOUT0#1	XI0/net1#3	1.14891e-18
C3057	XI0/XI1/Q#12	PHI#5	7.94002e-19
C3058	net7#19	SOUT1#11	9.00527e-19
C3059	net7#19	SOUT1#1	9.73491e-19
C3060	net7#17	SOUT1#6	1.79032e-18
C3061	SOUT1#22	net7#9	1.80819e-18
C3062	net7#2	SOUT1#3	2.27501e-18
C3063	VDD#144	SOUT2#20	5.92296e-19
C3064	VDD#62	SOUT2#6	6.94836e-19
C3065	SOUT2#11	VDD#149	7.64293e-19
C3066	SOUT2	VDD#113	7.94421e-19
C3067	VDD#68	SOUT2#1	1.21155e-18
C3068	SOUT2#11	VDD	1.24623e-18
C3069	SOUT2#8	VDD	2.30293e-18
C3070	VDD#152	SOUT2#1	2.33481e-18
C3071	XI0/XI1/D#14	SOUT0#4	7.99321e-19
C3072	XI0/XI1/D#2	SOUT0#4	8.55242e-19
C3073	XI0/XI1/D#15	SOUT0#5	1.40543e-18
C3074	VDD#133	SOUT3#20	5.92296e-19
C3075	VDD#88	SOUT3#6	6.94836e-19
C3076	SOUT3#11	VDD#138	7.64293e-19
C3077	SOUT3	VDD#106	7.94421e-19
C3078	VDD#94	SOUT3#1	1.21155e-18
C3079	SOUT3#11	VDD	1.24623e-18
C3080	SOUT3#8	VDD	2.30293e-18
C3081	VDD#141	SOUT3#1	2.33481e-18
C3082	XI3/XI0/XI1/net2#5	XI3/net1#10	3.92263e-19
C3083	XI0/XI0/XI0/BNOT#2	SOUT0#8	7.93386e-19
C3084	SOUT0#24	XI0/XI0/XI0/BNOT	8.11212e-19
C3085	XI0/XI0/XI0/BNOT#5	SOUT0#7	8.45903e-19
C3086	XI0/XI0/XI0/BNOT#10	SOUT0#3	9.04773e-19
C3087	SOUT0#22	XI0/XI0/XI0/BNOT#3	9.38469e-19
C3088	GND#64	net14#4	7.67752e-19
C3089	GND#46	net14#2	8.17588e-19
C3090	GND#99	net14#8	1.04902e-18
C3091	GND#137	net14#12	1.33266e-18
C3092	GND#50	net14#3	1.73249e-18
C3093	GND#66	net14#9	2.55369e-18
C3094	net7#5	VDD	5.05446e-19
C3095	VDD#50	net7#6	8.61141e-19
C3096	net7#21	VDD#26	1.06668e-18
C3097	net7#2	VDD#34	1.32554e-18
C3098	net7#19	VDD#161	1.41225e-18
C3099	VDD#166	net7#14	1.42169e-18
C3100	VDD#34	net7	1.73636e-18
C3101	net7#2	VDD	2.30792e-18
C3102	net7#2	VDD#27	2.42465e-18
C3103	VDD#165	net7	2.66145e-18
C3104	SOUT0#14	XI0/XI1/Q#2	9.16304e-19
C3105	XI1/XI1/D#15	GND#142	1.19132e-18
C3106	XI1/XI1/D#14	GND#141	1.22638e-18
C3107	XI2/XI1/D#12	XI2/net1#3	5.3688e-19
C3108	XI2/XI1/D#6	XI2/net1	5.92325e-19
C3109	XI2/XI1/D#16	XI2/net1	6.12214e-19
C3110	XI0/XI0/XI1/net2#13	SOUT0#4	4.31906e-19
C3111	XI0/XI0/XI1/net2#5	SOUT0#7	6.36383e-19
C3112	GND#34	XI1/XI1/XI4/net24#3	9.20398e-19
C3113	GND#34	XI1/XI1/XI4/net24#2	9.87977e-19
C3114	VDD#173	XI0/net1#4	7.43559e-19
C3115	VDD#172	XI0/net1#4	1.13006e-18
C3116	GND#106	XI1/XI0/XI0/BNOT#3	6.89259e-19
C3117	GND#106	XI1/XI0/XI0/BNOT#4	7.0191e-19
C3118	GND#138	XI1/XI1/Q#2	4.8289e-19
C3119	XI1/XI1/D#19	PHI#8	8.74572e-19
C3120	XI1/XI1/XI4/net24#2	PHI#12	7.75967e-19
C3121	XI1/XI1/XI4/net24#2	PHI#11	9.535e-19
C3122	XI0/XI0/XI0/BNOT#4	VDD#170	7.31422e-19
C3123	VDD#169	XI0/XI0/XI0/BNOT#3	1.12447e-18
C3124	XI0/XI0/XI0/BNOT#14	VDD#170	1.24021e-18
C3125	XI1/XI1/Q#12	PHI#11	7.94002e-19
C3126	XI3/XI1/D#20	XI3/XI1/Q	3.0256e-19
C3127	XI3/XI1/D#17	XI3/XI1/Q#3	3.77893e-19
C3128	XI3/XI1/Q#6	XI3/XI1/D#4	4.04483e-19
C3129	XI3/XI1/Q#5	XI3/XI1/D#3	4.90626e-19
C3130	XI3/XI1/D#17	XI3/XI1/Q#2	5.79029e-19
C3131	XI3/XI1/D#4	XI3/XI1/Q	6.8315e-19
C3132	XI0/XI1/D#12	XI0/net1#3	5.3688e-19
C3133	XI0/XI1/D#6	XI0/net1	5.92325e-19
C3134	XI0/XI1/D#16	XI0/net1	6.12214e-19
C3135	GND#86	net21#4	7.67752e-19
C3136	GND#68	net21#2	8.17588e-19
C3137	GND#92	net21#8	1.04902e-18
C3138	GND#128	net21#12	1.33266e-18
C3139	GND#72	net21#3	1.73249e-18
C3140	GND#88	net21#9	2.55369e-18
C3141	XI1/XI1/D#15	RST#6	1.25112e-18
C3142	XI2/XI1/D#15	GND#133	1.19132e-18
C3143	XI2/XI1/D#14	GND#132	1.22638e-18
C3144	GND#56	XI2/XI1/XI4/net24#3	9.20398e-19
C3145	GND#56	XI2/XI1/XI4/net24#2	9.87977e-19
C3146	GND#99	XI2/XI0/XI0/BNOT#3	6.89259e-19
C3147	GND#99	XI2/XI0/XI0/BNOT#4	7.0191e-19
C3148	VDD#166	XI0/XI0/XI1/net2#3	6.35307e-19
C3149	XI0/net1#16	XI0/XI0/XI0/BNOT#2	6.23458e-19
C3150	XI0/XI1/XI4/net24#12	XI0/XI1/XI4/PHINOT#2	5.31333e-19
C3151	COUT#5	XI3/XI0/XI1/net2	7.55169e-19
C3152	GND#129	XI2/XI1/Q#2	4.8289e-19
C3153	XI0/net1#16	XI0/XI0/XI0/ANOT#3	5.87684e-19
C3154	XI0/net1#6	XI0/XI0/XI0/ANOT	7.6486e-19
C3155	XI2/net1#16	XI2/XI0/XI0/BNOT#2	6.23458e-19
C3156	XI0/XI1/XI4/net24#4	XI0/XI1/D#4	6.43942e-19
C3157	XI0/XI1/XI4/net24#12	XI0/XI1/D#4	7.95905e-19
C3158	net7#14	XI0/XI0/XI1/net2	7.55169e-19
C3159	XI2/XI1/XI4/net24#12	XI2/XI1/XI4/PHINOT#2	5.31333e-19
C3160	SOUT1#2	XI1/net1#3	5.53224e-19
C3161	XI1/net1#2	SOUT1#1	5.64483e-19
C3162	XI1/net1#3	SOUT1#6	9.94394e-19
C3163	SOUT1#1	XI1/net1#3	1.14891e-18
C3164	XI0/XI0/XI1/net2#5	XI0/net1#10	3.92263e-19
C3165	XI2/XI1/D#19	PHI#14	8.74572e-19
C3166	XI3/XI1/XI4/net24#4	XI3/XI1/Q#2	6.00447e-19
C3167	XI3/XI0/XI0/BNOT#14	XI3/XI0/XI0/ANOT	6.36598e-19
C3168	XI3/XI0/XI0/BNOT#11	XI3/XI0/XI0/ANOT#2	7.40945e-19
C3169	XI2/XI1/XI4/net24#2	PHI#18	7.75967e-19
C3170	XI2/XI1/XI4/net24#2	PHI#17	9.535e-19
C3171	XI1/XI1/D#14	SOUT1#4	7.99321e-19
C3172	XI1/XI1/D#2	SOUT1#4	8.55242e-19
C3173	XI1/XI1/D#15	SOUT1#5	1.40543e-18
C3174	net14#19	SOUT2#11	9.00527e-19
C3175	net14#19	SOUT2#1	9.73491e-19
C3176	net14#17	SOUT2#6	1.79032e-18
C3177	SOUT2#22	net14#9	1.80819e-18
C3178	net14#2	SOUT2#3	2.27501e-18
C3179	XI3/XI1/D#15	GND#124	1.19132e-18
C3180	XI3/XI1/D#14	GND#123	1.22638e-18
C3181	XI2/XI1/Q#12	PHI#17	7.94002e-19
C3182	XI0/XI1/D#20	XI0/XI1/Q	3.0256e-19
C3183	XI0/XI1/D#17	XI0/XI1/Q#3	3.77893e-19
C3184	XI0/XI1/Q#6	XI0/XI1/D#4	4.04483e-19
C3185	XI0/XI1/Q#5	XI0/XI1/D#3	4.90626e-19
C3186	XI0/XI1/D#17	XI0/XI1/Q#2	5.79029e-19
C3187	XI0/XI1/D#4	XI0/XI1/Q	6.8315e-19
C3188	GND#78	XI3/XI1/XI4/net24#3	9.20398e-19
C3189	GND#78	XI3/XI1/XI4/net24#2	9.87977e-19
C3190	XI1/XI0/XI0/BNOT#2	SOUT1#8	7.93386e-19
C3191	SOUT1#24	XI1/XI0/XI0/BNOT	8.11212e-19
C3192	XI1/XI0/XI0/BNOT#5	SOUT1#7	8.45903e-19
C3193	XI1/XI0/XI0/BNOT#10	SOUT1#3	9.04773e-19
C3194	SOUT1#22	XI1/XI0/XI0/BNOT#3	9.38469e-19
C3195	XI2/net1#16	XI2/XI0/XI0/ANOT#3	5.87684e-19
C3196	XI2/net1#6	XI2/XI0/XI0/ANOT	7.6486e-19
C3197	GND#92	XI3/XI0/XI0/BNOT#3	6.89259e-19
C3198	GND#92	XI3/XI0/XI0/BNOT#4	7.03248e-19
C3199	XI2/XI1/XI4/net24#4	XI2/XI1/D#4	6.43942e-19
C3200	XI2/XI1/XI4/net24#12	XI2/XI1/D#4	7.95905e-19
C3201	XI2/net1#18	net14#9	3.7252e-19
C3202	XI2/net1#11	net14#6	3.75673e-19
C3203	XI2/net1#4	net14#17	4.08444e-19
C3204	XI2/net1#9	net14#7	7.33206e-19
C3205	XI2/net1#11	net14#7	7.62892e-19
C3206	XI2/net1#16	net14#9	9.2752e-19
C3207	GND#120	XI3/XI1/Q#2	4.8289e-19
C3208	XI0/XI1/XI4/net24#4	XI0/XI1/Q#2	6.00447e-19
C3209	SOUT1#14	XI1/XI1/Q#2	9.16304e-19
C3210	XI0/XI0/XI0/BNOT#14	XI0/XI0/XI0/ANOT	6.36598e-19
C3211	XI0/XI0/XI0/BNOT#11	XI0/XI0/XI0/ANOT#2	7.40945e-19
C3212	XI1/XI0/XI1/net2#13	SOUT1#4	4.31906e-19
C3213	XI1/XI0/XI1/net2#5	SOUT1#7	6.36383e-19
C3214	XI2/XI1/D#15	RST#9	1.25112e-18
C3215	net21#14	XI2/XI0/XI1/net2	7.55169e-19
C3216	net14#5	VDD	5.05446e-19
C3217	VDD#76	net14#6	8.61141e-19
C3218	net14#21	VDD#52	1.06668e-18
C3219	net14#2	VDD#60	1.32554e-18
C3220	net14#19	VDD#150	1.41225e-18
C3221	VDD#155	net14#14	1.42169e-18
C3222	VDD#60	net14	1.73636e-18
C3223	net14#2	VDD	2.30792e-18
C3224	net14#2	VDD#53	2.42465e-18
C3225	VDD#154	net14	2.66145e-18
C3226	VDD#162	XI1/net1#4	7.43559e-19
C3227	VDD#161	XI1/net1#4	1.13006e-18
C3228	XI3/XI1/D#19	PHI#20	8.74572e-19
C3229	XI2/XI1/D#14	net14#4	1.47002e-18
C3230	XI3/XI1/XI4/net24#2	PHI#24	7.75967e-19
C3231	XI3/XI1/XI4/net24#2	PHI#23	9.535e-19
C3232	XI3/XI1/Q#12	PHI#23	7.94002e-19
C3233	XI1/net1#18	net7#9	3.7252e-19
C3234	XI1/net1#11	net7#6	3.75673e-19
C3235	XI1/net1#4	net7#17	4.08444e-19
C3236	XI1/net1#9	net7#7	7.33206e-19
C3237	XI1/net1#11	net7#7	7.62892e-19
C3238	XI1/net1#16	net7#9	9.2752e-19
C3239	XI2/XI0/XI1/net2#5	XI2/net1#10	3.92263e-19
C3240	XI1/XI0/XI0/BNOT#4	VDD#159	7.31422e-19
C3241	VDD#158	XI1/XI0/XI0/BNOT#3	1.12447e-18
C3242	XI1/XI0/XI0/BNOT#14	VDD#159	1.24021e-18
C3243	XI1/XI1/D#14	net7#4	1.47002e-18
C3244	XI2/XI0/XI0/BNOT#5	net14	9.33843e-19
C3245	XI2/XI0/XI0/BNOT#7	net14#3	1.29331e-18
C3246	XI3/XI1/D#15	RST#12	1.25112e-18
C3247	VDD#155	XI1/XI0/XI1/net2#3	6.35307e-19
C3248	XI1/XI0/XI0/BNOT#5	net7	9.33843e-19
C3249	XI1/XI0/XI0/BNOT#7	net7#3	1.29331e-18
C3250	net7#19	XI1/XI0/XI0/ANOT	6.60017e-19
C3251	XI1/XI0/XI0/ANOT	net7#8	8.2626e-19
C3252	net14#19	XI2/XI0/XI0/ANOT	6.60017e-19
C3253	XI2/XI0/XI0/ANOT	net14#8	8.2626e-19
C3254	XI2/XI1/D#20	XI2/XI1/Q	3.0256e-19
C3255	XI2/XI1/D#17	XI2/XI1/Q#3	3.77893e-19
C3256	XI2/XI1/Q#6	XI2/XI1/D#4	4.04483e-19
C3257	XI2/XI1/Q#5	XI2/XI1/D#3	4.90626e-19
C3258	XI2/XI1/D#17	XI2/XI1/Q#2	5.79029e-19
C3259	XI2/XI1/D#4	XI2/XI1/Q	6.8315e-19
C3260	SOUT2#2	XI2/net1#3	5.53224e-19
C3261	XI2/net1#2	SOUT2#1	5.64483e-19
C3262	XI2/net1#3	SOUT2#6	9.94394e-19
C3263	SOUT2#1	XI2/net1#3	1.14891e-18
C3264	XI2/XI1/D#14	SOUT2#4	7.99321e-19
C3265	XI2/XI1/D#2	SOUT2#4	8.55242e-19
C3266	XI2/XI1/D#15	SOUT2#5	1.40543e-18
C3267	XI2/XI0/XI0/BNOT#2	SOUT2#8	7.93386e-19
C3268	SOUT2#24	XI2/XI0/XI0/BNOT	8.11212e-19
C3269	XI2/XI0/XI0/BNOT#5	SOUT2#7	8.45903e-19
C3270	XI2/XI0/XI0/BNOT#10	SOUT2#3	9.04773e-19
C3271	SOUT2#22	XI2/XI0/XI0/BNOT#3	9.38469e-19
C3272	net21#19	SOUT3#11	9.00527e-19
C3273	net21#19	SOUT3#1	9.73491e-19
C3274	net21#17	SOUT3#6	1.79032e-18
C3275	SOUT3#22	net21#9	1.80819e-18
C3276	net21#2	SOUT3#3	2.27501e-18
C3277	XI2/XI1/XI4/net24#4	XI2/XI1/Q#2	6.00447e-19
C3278	SOUT2#14	XI2/XI1/Q#2	9.16304e-19
C3279	XI2/XI0/XI0/BNOT#14	XI2/XI0/XI0/ANOT	6.36598e-19
C3280	XI2/XI0/XI0/BNOT#11	XI2/XI0/XI0/ANOT#2	7.40945e-19
C3281	XI2/XI0/XI1/net2#13	SOUT2#4	4.31906e-19
C3282	XI2/XI0/XI1/net2#5	SOUT2#7	6.36383e-19
C3283	net21#5	VDD	5.05446e-19
C3284	VDD#102	net21#6	8.61141e-19
C3285	net21#21	VDD#78	1.06668e-18
C3286	net21#2	VDD#86	1.32554e-18
C3287	net21#19	VDD#139	1.41225e-18
C3288	VDD#144	net21#14	1.42169e-18
C3289	VDD#86	net21	1.73636e-18
C3290	net21#2	VDD	2.30792e-18
C3291	net21#2	VDD#79	2.42465e-18
C3292	VDD#143	net21	2.66145e-18
C3293	VDD#151	XI2/net1#4	7.43559e-19
C3294	VDD#150	XI2/net1#4	1.13006e-18
C3295	XI2/XI0/XI0/BNOT#4	VDD#148	7.31422e-19
C3296	VDD#147	XI2/XI0/XI0/BNOT#3	1.12447e-18
C3297	XI2/XI0/XI0/BNOT#14	VDD#148	1.24021e-18
C3298	VDD#144	XI2/XI0/XI1/net2#3	6.35307e-19
C3299	SOUT3#2	XI3/net1#3	5.53224e-19
C3300	XI3/net1#2	SOUT3#1	5.64483e-19
C3301	XI3/net1#3	SOUT3#6	9.94394e-19
C3302	SOUT3#1	XI3/net1#3	1.14891e-18
C3303	XI3/XI1/D#14	SOUT3#4	7.99321e-19
C3304	XI3/XI1/D#2	SOUT3#4	8.55242e-19
C3305	XI3/XI1/D#15	SOUT3#5	1.40543e-18
C3306	XI3/XI0/XI0/BNOT#2	SOUT3#8	7.93386e-19
C3307	SOUT3#24	XI3/XI0/XI0/BNOT	8.11212e-19
C3308	XI3/XI0/XI0/BNOT#5	SOUT3#7	8.45903e-19
C3309	XI3/XI0/XI0/BNOT#10	SOUT3#3	9.04773e-19
C3310	SOUT3#22	XI3/XI0/XI0/BNOT#3	9.38469e-19
C3311	SOUT3#14	XI3/XI1/Q#2	9.16304e-19
C3312	VDD#140	XI3/net1#4	7.43559e-19
C3313	VDD#139	XI3/net1#4	1.13006e-18
C3314	XI3/XI0/XI1/net2#13	SOUT3#4	4.31906e-19
C3315	XI3/XI0/XI1/net2#5	SOUT3#7	6.36383e-19
C3316	XI3/XI0/XI0/BNOT#4	VDD#137	7.31422e-19
C3317	VDD#136	XI3/XI0/XI0/BNOT#3	1.12447e-18
C3318	XI3/XI0/XI0/BNOT#14	VDD#137	1.24021e-18
C3319	VDD#133	XI3/XI0/XI1/net2#3	6.35307e-19
C3320	XI3/net1#18	net21#9	3.7252e-19
C3321	XI3/net1#11	net21#6	3.75673e-19
C3322	XI3/net1#4	net21#17	4.08444e-19
C3323	XI3/net1#9	net21#7	7.33206e-19
C3324	XI3/net1#11	net21#7	7.62892e-19
C3325	XI3/net1#16	net21#9	9.2752e-19
C3326	XI3/XI1/D#14	net21#4	1.47002e-18
C3327	XI3/XI1/D#12	XI3/net1#3	5.3688e-19
C3328	XI3/XI1/D#6	XI3/net1	5.92325e-19
C3329	XI3/XI1/D#16	XI3/net1	6.12214e-19
C3330	XI3/XI0/XI0/BNOT#5	net21	9.33843e-19
C3331	XI3/XI0/XI0/BNOT#7	net21#3	1.29331e-18
C3332	XI1/XI1/D#12	XI1/net1#3	5.3688e-19
C3333	XI1/XI1/D#6	XI1/net1	5.92325e-19
C3334	XI1/XI1/D#16	XI1/net1	6.12214e-19
C3335	net21#19	XI3/XI0/XI0/ANOT	6.60017e-19
C3336	XI3/XI0/XI0/ANOT	net21#8	8.2626e-19
C3337	XI1/net1#16	XI1/XI0/XI0/BNOT#2	6.23458e-19
C3338	XI1/XI1/XI4/net24#12	XI1/XI1/XI4/PHINOT#2	5.31333e-19
C3339	XI1/net1#16	XI1/XI0/XI0/ANOT#3	5.87684e-19
C3340	XI1/net1#6	XI1/XI0/XI0/ANOT	7.6486e-19
C3341	XI3/net1#16	XI3/XI0/XI0/BNOT#2	6.23458e-19
C3342	XI1/XI1/XI4/net24#4	XI1/XI1/D#4	6.43942e-19
C3343	XI1/XI1/XI4/net24#12	XI1/XI1/D#4	7.95905e-19
C3344	XI3/XI1/XI4/net24#12	XI3/XI1/XI4/PHINOT#2	5.31333e-19
C3345	net14#14	XI1/XI0/XI1/net2	7.55169e-19
C3346	XI1/XI0/XI1/net2#5	XI1/net1#10	3.92263e-19
C3347	XI3/net1#16	XI3/XI0/XI0/ANOT#3	5.87684e-19
C3348	XI3/net1#6	XI3/XI0/XI0/ANOT	7.6486e-19
C3349	XI3/XI1/XI4/net24#4	XI3/XI1/D#4	6.43942e-19
C3350	XI3/XI1/XI4/net24#12	XI3/XI1/D#4	7.95905e-19
C3351	CIN	GND	5.37703e-17
C3352	COUT	GND	7.19493e-17
C3353	PHI	GND	3.10368e-17
C3354	RST	GND	4.28879e-17
C3355	SOUT0	GND	1.90083e-17
C3356	SOUT1	GND	1.90083e-17
C3357	SOUT2	GND	1.90083e-17
C3358	SOUT3	GND	1.90083e-17
C3359	VDD	GND	2.52104e-18
C3360	XI0/XI0/XI0/net4	GND	3.66456e-19
C3361	XI0/XI1/XI4/net9	GND	3.18655e-19
C3362	XI0/XI1/XI4/net25	GND	3.17892e-19
C3363	XI1/XI0/XI0/net4	GND	3.66456e-19
C3364	XI1/XI1/XI4/net9	GND	3.18655e-19
C3365	XI1/XI1/XI4/net25	GND	3.17892e-19
C3366	XI2/XI0/XI0/net4	GND	3.66456e-19
C3367	XI2/XI1/XI4/net9	GND	3.18655e-19
C3368	XI2/XI1/XI4/net25	GND	3.17892e-19
C3369	XI3/XI0/XI0/net4	GND	3.66456e-19
C3370	XI3/XI1/XI4/net9	GND	3.18655e-19
C3371	XI3/XI1/XI4/net25	GND	3.17892e-19
C3372	XI3/XI0/XI1/net2#3	GND	3.13736e-18
C3373	XI3/XI0/XI0/BNOT#3	GND	1.96891e-18
C3374	XI3/XI1/Q	GND	2.6773e-18
C3375	net21#7	GND	4.03466e-18
C3376	PHI#22	GND	1.97867e-18
C3377	XI3/XI1/D#3	GND	2.28632e-20
C3378	net21#6	GND	1.53502e-18
C3379	XI3/XI0/XI0/ANOT	GND	1.42922e-17
C3380	SOUT3#7	GND	6.82093e-19
C3381	XI3/XI1/XI4/net24	GND	4.03648e-18
C3382	XI3/XI1/XI4/PHINOT	GND	4.28642e-19
C3383	SOUT3#6	GND	7.98051e-18
C3384	XI3/net1#3	GND	1.99398e-18
C3385	SOUT3#1	GND	5.3701e-19
C3386	RST#12	GND	2.45689e-17
C3387	net21	GND	2.83442e-18
C3388	XI2/XI0/XI1/net2#3	GND	3.13736e-18
C3389	XI2/XI0/XI0/BNOT#3	GND	1.96891e-18
C3390	XI2/XI1/Q	GND	2.6773e-18
C3391	net14#7	GND	4.03466e-18
C3392	PHI#16	GND	1.97867e-18
C3393	XI2/XI1/D#3	GND	2.28632e-20
C3394	net14#6	GND	1.53502e-18
C3395	XI2/XI0/XI0/ANOT	GND	1.42922e-17
C3396	SOUT2#7	GND	6.82093e-19
C3397	XI2/XI1/XI4/net24	GND	4.03648e-18
C3398	XI2/XI1/XI4/PHINOT	GND	4.28642e-19
C3399	SOUT2#6	GND	7.98051e-18
C3400	XI2/net1#3	GND	1.99398e-18
C3401	SOUT2#1	GND	5.3701e-19
C3402	RST#9	GND	2.45689e-17
C3403	net14	GND	2.83442e-18
C3404	XI1/XI0/XI1/net2#3	GND	3.13736e-18
C3405	XI1/XI0/XI0/BNOT#3	GND	1.96891e-18
C3406	XI1/XI1/Q	GND	2.6773e-18
C3407	net7#7	GND	4.03466e-18
C3408	PHI#10	GND	1.97867e-18
C3409	XI1/XI1/D#3	GND	2.28632e-20
C3410	net7#6	GND	1.53502e-18
C3411	XI1/XI0/XI0/ANOT	GND	1.42922e-17
C3412	SOUT1#7	GND	6.82093e-19
C3413	XI1/XI1/XI4/net24	GND	4.03648e-18
C3414	XI1/XI1/XI4/PHINOT	GND	4.28642e-19
C3415	SOUT1#6	GND	7.98051e-18
C3416	XI1/net1#3	GND	1.99398e-18
C3417	SOUT1#1	GND	5.3701e-19
C3418	RST#6	GND	2.45689e-17
C3419	net7	GND	2.83442e-18
C3420	XI0/XI0/XI1/net2#3	GND	3.13736e-18
C3421	XI0/XI0/XI0/BNOT#3	GND	1.96891e-18
C3422	XI0/XI1/Q	GND	2.6773e-18
C3423	CIN#7	GND	4.03466e-18
C3424	PHI#4	GND	1.97867e-18
C3425	XI0/XI1/D#3	GND	2.28632e-20
C3426	CIN#6	GND	1.05456e-18
C3427	XI0/XI0/XI0/ANOT	GND	1.42922e-17
C3428	SOUT0#7	GND	6.82093e-19
C3429	XI0/XI1/XI4/net24	GND	4.03648e-18
C3430	XI0/XI1/XI4/PHINOT	GND	4.28642e-19
C3431	SOUT0#6	GND	7.98051e-18
C3432	XI0/net1#3	GND	1.99398e-18
C3433	SOUT0#1	GND	5.3701e-19
C3434	RST#3	GND	2.33004e-17
C3435	CIN#1	GND	2.83442e-18
C3436	XI3/XI0/XI1/net2	GND	2.79716e-17
C3437	SOUT3#9	GND	6.61416e-18
C3438	XI3/XI1/Q#3	GND	1.48647e-17
C3439	net21#9	GND	1.32586e-17
C3440	PHI#24	GND	2.01904e-17
C3441	XI3/XI1/XI4/net24#3	GND	9.99763e-18
C3442	net21#4	GND	3.26818e-17
C3443	XI3/XI0/XI0/ANOT#3	GND	1.01721e-17
C3444	XI3/XI0/XI0/BNOT	GND	6.49394e-18
C3445	XI3/XI1/D	GND	6.5331e-18
C3446	XI3/XI1/XI4/PHINOT#3	GND	1.96485e-17
C3447	SOUT3#4	GND	1.86891e-17
C3448	XI3/net1	GND	3.35095e-17
C3449	SOUT3#3	GND	2.75159e-17
C3450	PHI#21	GND	5.87414e-17
C3451	RST#10	GND	1.1724e-17
C3452	net21#3	GND	3.0384e-17
C3453	XI2/XI0/XI1/net2	GND	3.01059e-17
C3454	SOUT2#9	GND	6.61416e-18
C3455	XI2/XI1/Q#3	GND	1.48647e-17
C3456	net14#9	GND	1.32586e-17
C3457	PHI#18	GND	1.88184e-17
C3458	XI2/XI1/XI4/net24#3	GND	9.99763e-18
C3459	net14#4	GND	3.26818e-17
C3460	XI2/XI0/XI0/ANOT#3	GND	1.01721e-17
C3461	XI2/XI0/XI0/BNOT	GND	6.49394e-18
C3462	XI2/XI1/D	GND	6.5331e-18
C3463	XI2/XI1/XI4/PHINOT#3	GND	1.96485e-17
C3464	SOUT2#4	GND	1.86891e-17
C3465	XI2/net1	GND	3.35095e-17
C3466	SOUT2#3	GND	2.75159e-17
C3467	PHI#15	GND	5.87414e-17
C3468	RST#7	GND	1.1724e-17
C3469	net14#3	GND	3.0384e-17
C3470	XI1/XI0/XI1/net2	GND	3.01059e-17
C3471	SOUT1#9	GND	6.61416e-18
C3472	XI1/XI1/Q#3	GND	1.48647e-17
C3473	net7#9	GND	1.32586e-17
C3474	PHI#12	GND	1.88184e-17
C3475	XI1/XI1/XI4/net24#3	GND	9.99763e-18
C3476	net7#4	GND	3.26818e-17
C3477	XI1/XI0/XI0/ANOT#3	GND	1.01721e-17
C3478	XI1/XI0/XI0/BNOT	GND	6.49394e-18
C3479	XI1/XI1/D	GND	6.5331e-18
C3480	XI1/XI1/XI4/PHINOT#3	GND	1.96485e-17
C3481	SOUT1#4	GND	1.86891e-17
C3482	XI1/net1	GND	3.35095e-17
C3483	SOUT1#3	GND	2.75159e-17
C3484	PHI#9	GND	5.87414e-17
C3485	RST#4	GND	1.1724e-17
C3486	net7#3	GND	3.0384e-17
C3487	XI0/XI0/XI1/net2	GND	3.01059e-17
C3488	SOUT0#9	GND	6.61416e-18
C3489	XI0/XI1/Q#3	GND	1.48647e-17
C3490	CIN#9	GND	1.2684e-17
C3491	PHI#6	GND	1.88184e-17
C3492	XI0/XI1/XI4/net24#3	GND	9.99763e-18
C3493	CIN#4	GND	3.26818e-17
C3494	XI0/XI0/XI0/ANOT#3	GND	1.01721e-17
C3495	XI0/XI0/XI0/BNOT	GND	6.49394e-18
C3496	XI0/XI1/D	GND	6.5331e-18
C3497	XI0/XI1/XI4/PHINOT#3	GND	1.96485e-17
C3498	SOUT0#4	GND	1.86891e-17
C3499	XI0/net1	GND	3.35095e-17
C3500	SOUT0#3	GND	2.75159e-17
C3501	PHI#3	GND	5.87414e-17
C3502	RST#1	GND	1.1724e-17
C3503	CIN#3	GND	3.0384e-17
C3504	XI3/XI0/XI0/BNOT#4	GND	1.36471e-17
C3505	SOUT3#10	GND	2.91212e-17
C3506	XI3/XI0/XI1/net2#2	GND	4.81417e-17
C3507	XI3/XI1/Q#2	GND	5.16577e-17
C3508	net21#8	GND	5.85133e-17
C3509	PHI#23	GND	5.15321e-17
C3510	XI3/XI1/D#4	GND	4.17494e-19
C3511	XI3/XI1/XI4/net24#4	GND	1.30667e-17
C3512	net21#5	GND	4.82674e-17
C3513	XI3/XI0/XI0/ANOT#2	GND	7.68838e-17
C3514	SOUT3#8	GND	2.47258e-17
C3515	XI3/XI0/XI0/BNOT#2	GND	2.18423e-17
C3516	XI3/XI1/XI4/net24#2	GND	1.89551e-17
C3517	XI3/XI1/D#2	GND	1.32495e-17
C3518	XI3/XI1/XI4/PHINOT#2	GND	5.17685e-17
C3519	SOUT3#5	GND	7.09963e-17
C3520	XI3/net1#2	GND	2.87717e-17
C3521	SOUT3#2	GND	4.38104e-17
C3522	PHI#20	GND	1.18812e-16
C3523	RST#11	GND	2.11303e-16
C3524	net21#2	GND	1.38027e-16
C3525	XI2/XI0/XI0/BNOT#4	GND	1.36298e-17
C3526	SOUT2#10	GND	2.91212e-17
C3527	XI2/XI0/XI1/net2#2	GND	4.81417e-17
C3528	XI2/XI1/Q#2	GND	5.16577e-17
C3529	net14#8	GND	5.85174e-17
C3530	PHI#17	GND	6.63162e-17
C3531	XI2/XI1/D#4	GND	4.17494e-19
C3532	XI2/XI1/XI4/net24#4	GND	1.30667e-17
C3533	net14#5	GND	4.82674e-17
C3534	XI2/XI0/XI0/ANOT#2	GND	7.68838e-17
C3535	SOUT2#8	GND	2.47258e-17
C3536	XI2/XI0/XI0/BNOT#2	GND	2.18423e-17
C3537	XI2/XI1/XI4/net24#2	GND	1.89551e-17
C3538	XI2/XI1/D#2	GND	1.32495e-17
C3539	XI2/XI1/XI4/PHINOT#2	GND	5.17685e-17
C3540	SOUT2#5	GND	7.03277e-17
C3541	XI2/net1#2	GND	2.87717e-17
C3542	SOUT2#2	GND	4.38104e-17
C3543	PHI#14	GND	1.18812e-16
C3544	RST#8	GND	2.24025e-16
C3545	net14#2	GND	1.38027e-16
C3546	XI1/XI0/XI0/BNOT#4	GND	1.36298e-17
C3547	SOUT1#10	GND	2.91212e-17
C3548	XI1/XI0/XI1/net2#2	GND	4.81417e-17
C3549	XI1/XI1/Q#2	GND	5.16577e-17
C3550	net7#8	GND	5.85174e-17
C3551	PHI#11	GND	6.63162e-17
C3552	XI1/XI1/D#4	GND	4.17494e-19
C3553	XI1/XI1/XI4/net24#4	GND	1.30667e-17
C3554	net7#5	GND	4.82674e-17
C3555	XI1/XI0/XI0/ANOT#2	GND	7.68838e-17
C3556	SOUT1#8	GND	2.47258e-17
C3557	XI1/XI0/XI0/BNOT#2	GND	2.18423e-17
C3558	XI1/XI1/XI4/net24#2	GND	1.89551e-17
C3559	XI1/XI1/D#2	GND	1.32495e-17
C3560	XI1/XI1/XI4/PHINOT#2	GND	5.17685e-17
C3561	SOUT1#5	GND	7.03277e-17
C3562	XI1/net1#2	GND	2.87717e-17
C3563	SOUT1#2	GND	4.38104e-17
C3564	PHI#8	GND	1.18812e-16
C3565	RST#5	GND	2.24025e-16
C3566	net7#2	GND	1.38027e-16
C3567	XI0/XI0/XI0/BNOT#4	GND	1.36298e-17
C3568	SOUT0#10	GND	2.91212e-17
C3569	XI0/XI0/XI1/net2#2	GND	4.81417e-17
C3570	XI0/XI1/Q#2	GND	5.16577e-17
C3571	CIN#8	GND	5.85367e-17
C3572	PHI#5	GND	6.63162e-17
C3573	XI0/XI1/D#4	GND	4.17494e-19
C3574	XI0/XI1/XI4/net24#4	GND	1.30667e-17
C3575	CIN#5	GND	4.82674e-17
C3576	XI0/XI0/XI0/ANOT#2	GND	7.68838e-17
C3577	SOUT0#8	GND	2.47258e-17
C3578	XI0/XI0/XI0/BNOT#2	GND	2.18423e-17
C3579	XI0/XI1/XI4/net24#2	GND	1.89551e-17
C3580	XI0/XI1/D#2	GND	1.32495e-17
C3581	XI0/XI1/XI4/PHINOT#2	GND	5.17685e-17
C3582	SOUT0#5	GND	7.03277e-17
C3583	XI0/net1#2	GND	2.87717e-17
C3584	SOUT0#2	GND	4.38104e-17
C3585	PHI#2	GND	6.66514e-17
C3586	RST#2	GND	1.17958e-16
C3587	CIN#2	GND	8.12975e-17
C3588	VDD#105	GND	6.12471e-17
C3589	VDD#133	GND	5.19488e-17
C3590	COUT#5	GND	2.8667e-17
C3591	COUT#7	GND	4.17009e-17
C3592	SOUT3#18	GND	4.38955e-17
C3593	SOUT3#20	GND	6.34514e-17
C3594	SOUT3#22	GND	3.17463e-17
C3595	COUT#3	GND	8.67498e-18
C3596	COUT#6	GND	1.18863e-17
C3597	COUT#1	GND	1.10923e-17
C3598	SOUT3#14	GND	3.23603e-18
C3599	SOUT3#19	GND	1.94159e-17
C3600	SOUT3#16	GND	8.43156e-18
C3601	VDD#104	GND	3.11409e-18
C3602	VDD#102	GND	2.60645e-19
C3603	VDD#137	GND	2.30328e-19
C3604	VDD#100	GND	2.25295e-18
C3605	XI3/net1#6	GND	3.57652e-19
C3606	XI3/XI0/XI0/BNOT#14	GND	9.80305e-18
C3607	XI3/XI0/XI0/BNOT#9	GND	3.05937e-17
C3608	XI3/XI0/XI0/BNOT#11	GND	1.8348e-17
C3609	XI3/XI0/XI1/net2#13	GND	1.75343e-17
C3610	XI3/XI0/XI1/net2#15	GND	2.92719e-17
C3611	XI3/net1#4	GND	6.20306e-18
C3612	XI3/net1#9	GND	7.68836e-18
C3613	XI3/net1#16	GND	2.01534e-17
C3614	XI3/XI1/XI4/net24#11	GND	2.17241e-18
C3615	XI3/XI1/XI4/net24#12	GND	1.17061e-17
C3616	XI3/XI1/Q#11	GND	2.17936e-17
C3617	XI3/XI1/Q#9	GND	1.09498e-17
C3618	XI3/XI0/XI1/net2#12	GND	8.07284e-18
C3619	VDD#98	GND	3.74949e-19
C3620	VDD#138	GND	3.8563e-19
C3621	VDD#96	GND	1.60408e-18
C3622	SOUT3#11	GND	1.47001e-17
C3623	SOUT3#24	GND	1.94621e-17
C3624	XI3/XI1/D#20	GND	3.08439e-18
C3625	XI3/XI1/D#17	GND	1.03658e-17
C3626	XI3/XI0/XI1/net2#16	GND	6.12784e-18
C3627	XI3/XI1/Q#6	GND	4.30485e-18
C3628	XI3/XI1/Q#12	GND	1.07738e-17
C3629	VDD#139	GND	2.20938e-19
C3630	VDD#94	GND	1.74327e-18
C3631	VDD#110	GND	2.81797e-20
C3632	VDD#92	GND	6.91838e-19
C3633	XI3/XI0/XI1/XI0/net13#4	GND	1.30885e-17
C3634	XI3/XI0/XI1/net2#9	GND	6.73319e-19
C3635	XI3/XI1/Q#5	GND	2.09121e-18
C3636	XI3/XI1/Q#7	GND	2.16707e-19
C3637	XI3/XI1/XI4/net24#13	GND	1.93822e-17
C3638	XI3/XI1/XI4/net24#6	GND	7.33241e-18
C3639	XI3/XI1/XI4/net24#9	GND	1.65682e-17
C3640	VDD#90	GND	1.17069e-18
C3641	XI3/XI1/D#19	GND	3.36909e-17
C3642	XI3/XI1/D#14	GND	2.50795e-17
C3643	net21#17	GND	2.67287e-17
C3644	net21#19	GND	4.2371e-17
C3645	VDD#88	GND	4.14886e-19
C3646	XI3/XI0/XI0/BNOT#5	GND	1.84278e-19
C3647	XI3/XI0/XI0/BNOT#10	GND	3.17641e-17
C3648	XI3/XI0/XI0/BNOT#7	GND	2.10842e-17
C3649	XI3/XI1/D#7	GND	8.64157e-19
C3650	XI3/XI1/XI5/net13#3	GND	1.06358e-17
C3651	VDD#142	GND	1.23331e-18
C3652	VDD#86	GND	2.68286e-19
C3653	XI3/XI1/D#15	GND	3.82381e-17
C3654	XI3/XI1/D#10	GND	6.97924e-18
C3655	XI3/XI1/XI4/PHINOT#4	GND	1.77609e-18
C3656	XI3/XI1/XI4/PHINOT#9	GND	5.23298e-17
C3657	XI3/XI1/XI4/PHINOT#6	GND	2.42089e-17
C3658	XI3/XI0/XI0/ANOT#4	GND	9.81082e-18
C3659	XI3/XI0/XI0/ANOT#9	GND	4.88348e-17
C3660	XI3/XI0/XI0/ANOT#6	GND	1.02907e-17
C3661	VDD#83	GND	3.60805e-19
C3662	VDD#82	GND	1.26825e-18
C3663	XI3/XI1/D#6	GND	1.74398e-17
C3664	XI3/XI1/D#16	GND	2.45897e-17
C3665	VDD#143	GND	7.14874e-20
C3666	VDD#80	GND	8.37146e-19
C3667	VDD#112	GND	5.95395e-17
C3668	VDD#144	GND	4.90747e-17
C3669	net21#14	GND	2.8667e-17
C3670	net21#21	GND	8.96238e-17
C3671	SOUT2#18	GND	4.38955e-17
C3672	SOUT2#20	GND	6.30224e-17
C3673	SOUT2#22	GND	3.18348e-17
C3674	net21#12	GND	8.67498e-18
C3675	net21#15	GND	1.18863e-17
C3676	net21#10	GND	1.10923e-17
C3677	SOUT2#14	GND	3.23603e-18
C3678	SOUT2#19	GND	1.94159e-17
C3679	SOUT2#16	GND	8.43156e-18
C3680	VDD#78	GND	3.11409e-18
C3681	VDD#76	GND	2.60645e-19
C3682	VDD#148	GND	2.30328e-19
C3683	VDD#74	GND	2.25295e-18
C3684	XI2/net1#6	GND	3.57652e-19
C3685	XI2/XI0/XI0/BNOT#14	GND	9.80305e-18
C3686	XI2/XI0/XI0/BNOT#9	GND	3.07644e-17
C3687	XI2/XI0/XI0/BNOT#11	GND	1.8348e-17
C3688	XI2/XI0/XI1/net2#13	GND	1.75343e-17
C3689	XI2/XI0/XI1/net2#15	GND	2.92719e-17
C3690	XI2/net1#4	GND	6.20306e-18
C3691	XI2/net1#9	GND	7.68836e-18
C3692	XI2/net1#16	GND	2.01534e-17
C3693	XI2/XI1/XI4/net24#11	GND	2.17241e-18
C3694	XI2/XI1/XI4/net24#12	GND	1.17061e-17
C3695	XI2/XI1/Q#11	GND	2.17936e-17
C3696	XI2/XI1/Q#9	GND	1.09498e-17
C3697	XI2/XI0/XI1/net2#12	GND	8.07284e-18
C3698	VDD#72	GND	3.74949e-19
C3699	VDD#149	GND	3.8563e-19
C3700	VDD#70	GND	1.60408e-18
C3701	SOUT2#11	GND	1.47001e-17
C3702	SOUT2#24	GND	1.94621e-17
C3703	XI2/XI1/D#20	GND	3.08439e-18
C3704	XI2/XI1/D#17	GND	1.03658e-17
C3705	XI2/XI0/XI1/net2#16	GND	6.12784e-18
C3706	XI2/XI1/Q#6	GND	4.30485e-18
C3707	XI2/XI1/Q#12	GND	1.07738e-17
C3708	VDD#150	GND	2.20938e-19
C3709	VDD#68	GND	1.74327e-18
C3710	VDD#117	GND	2.81797e-20
C3711	VDD#66	GND	6.91838e-19
C3712	XI2/XI0/XI1/XI0/net13#4	GND	1.30885e-17
C3713	XI2/XI0/XI1/net2#9	GND	6.73319e-19
C3714	XI2/XI1/Q#5	GND	2.09121e-18
C3715	XI2/XI1/Q#7	GND	2.16707e-19
C3716	XI2/XI1/XI4/net24#13	GND	1.93822e-17
C3717	XI2/XI1/XI4/net24#6	GND	7.33241e-18
C3718	XI2/XI1/XI4/net24#9	GND	1.65682e-17
C3719	VDD#64	GND	1.17069e-18
C3720	XI2/XI1/D#19	GND	3.36909e-17
C3721	XI2/XI1/D#14	GND	2.50795e-17
C3722	net14#17	GND	2.67287e-17
C3723	net14#19	GND	4.2371e-17
C3724	VDD#62	GND	4.14886e-19
C3725	XI2/XI0/XI0/BNOT#5	GND	1.84278e-19
C3726	XI2/XI0/XI0/BNOT#10	GND	3.17641e-17
C3727	XI2/XI0/XI0/BNOT#7	GND	2.10842e-17
C3728	XI2/XI1/D#7	GND	8.64157e-19
C3729	XI2/XI1/XI5/net13#3	GND	1.06358e-17
C3730	VDD#153	GND	1.23331e-18
C3731	VDD#60	GND	2.68286e-19
C3732	XI2/XI1/D#15	GND	3.82381e-17
C3733	XI2/XI1/D#10	GND	6.97924e-18
C3734	XI2/XI1/XI4/PHINOT#4	GND	1.77609e-18
C3735	XI2/XI1/XI4/PHINOT#9	GND	5.23298e-17
C3736	XI2/XI1/XI4/PHINOT#6	GND	2.42089e-17
C3737	XI2/XI0/XI0/ANOT#4	GND	9.81082e-18
C3738	XI2/XI0/XI0/ANOT#9	GND	4.88348e-17
C3739	XI2/XI0/XI0/ANOT#6	GND	1.02907e-17
C3740	VDD#57	GND	3.60805e-19
C3741	VDD#56	GND	1.26825e-18
C3742	XI2/XI1/D#6	GND	1.74398e-17
C3743	XI2/XI1/D#16	GND	2.45897e-17
C3744	VDD#154	GND	7.14874e-20
C3745	VDD#54	GND	8.37146e-19
C3746	VDD#119	GND	5.95395e-17
C3747	VDD#155	GND	4.90747e-17
C3748	net14#14	GND	2.8667e-17
C3749	net14#21	GND	8.96238e-17
C3750	SOUT1#18	GND	4.38955e-17
C3751	SOUT1#20	GND	6.30224e-17
C3752	SOUT1#22	GND	3.18348e-17
C3753	net14#12	GND	8.67498e-18
C3754	net14#15	GND	1.18863e-17
C3755	net14#10	GND	1.10923e-17
C3756	SOUT1#14	GND	3.23603e-18
C3757	SOUT1#19	GND	1.94159e-17
C3758	SOUT1#16	GND	8.43156e-18
C3759	VDD#52	GND	3.11409e-18
C3760	VDD#50	GND	2.60645e-19
C3761	VDD#159	GND	2.30328e-19
C3762	VDD#48	GND	2.25295e-18
C3763	XI1/net1#6	GND	3.57652e-19
C3764	XI1/XI0/XI0/BNOT#14	GND	9.80305e-18
C3765	XI1/XI0/XI0/BNOT#9	GND	3.07644e-17
C3766	XI1/XI0/XI0/BNOT#11	GND	1.8348e-17
C3767	XI1/XI0/XI1/net2#13	GND	1.75343e-17
C3768	XI1/XI0/XI1/net2#15	GND	2.92719e-17
C3769	XI1/net1#4	GND	6.20306e-18
C3770	XI1/net1#9	GND	7.68836e-18
C3771	XI1/net1#16	GND	2.01534e-17
C3772	XI1/XI1/XI4/net24#11	GND	2.17241e-18
C3773	XI1/XI1/XI4/net24#12	GND	1.17061e-17
C3774	XI1/XI1/Q#11	GND	2.17936e-17
C3775	XI1/XI1/Q#9	GND	1.09498e-17
C3776	XI1/XI0/XI1/net2#12	GND	8.07284e-18
C3777	VDD#46	GND	3.74949e-19
C3778	VDD#160	GND	3.8563e-19
C3779	VDD#44	GND	1.60408e-18
C3780	SOUT1#11	GND	1.47001e-17
C3781	SOUT1#24	GND	1.94621e-17
C3782	XI1/XI1/D#20	GND	3.08439e-18
C3783	XI1/XI1/D#17	GND	1.03658e-17
C3784	XI1/XI0/XI1/net2#16	GND	6.12784e-18
C3785	XI1/XI1/Q#6	GND	4.30485e-18
C3786	XI1/XI1/Q#12	GND	1.07738e-17
C3787	VDD#161	GND	2.20938e-19
C3788	VDD#42	GND	1.74327e-18
C3789	VDD#124	GND	2.81797e-20
C3790	VDD#40	GND	6.91838e-19
C3791	XI1/XI0/XI1/XI0/net13#4	GND	1.30885e-17
C3792	XI1/XI0/XI1/net2#9	GND	6.73319e-19
C3793	XI1/XI1/Q#5	GND	2.09121e-18
C3794	XI1/XI1/Q#7	GND	2.16707e-19
C3795	XI1/XI1/XI4/net24#13	GND	1.93822e-17
C3796	XI1/XI1/XI4/net24#6	GND	7.33241e-18
C3797	XI1/XI1/XI4/net24#9	GND	1.65682e-17
C3798	VDD#38	GND	1.17069e-18
C3799	XI1/XI1/D#19	GND	3.36909e-17
C3800	XI1/XI1/D#14	GND	2.50795e-17
C3801	net7#17	GND	2.67287e-17
C3802	net7#19	GND	4.2371e-17
C3803	VDD#36	GND	4.14886e-19
C3804	XI1/XI0/XI0/BNOT#5	GND	1.84278e-19
C3805	XI1/XI0/XI0/BNOT#10	GND	3.17641e-17
C3806	XI1/XI0/XI0/BNOT#7	GND	2.10842e-17
C3807	XI1/XI1/D#7	GND	8.64157e-19
C3808	XI1/XI1/XI5/net13#3	GND	1.06358e-17
C3809	VDD#164	GND	1.23331e-18
C3810	VDD#34	GND	2.68286e-19
C3811	XI1/XI1/D#15	GND	3.82381e-17
C3812	XI1/XI1/D#10	GND	6.97924e-18
C3813	XI1/XI1/XI4/PHINOT#4	GND	1.77609e-18
C3814	XI1/XI1/XI4/PHINOT#9	GND	5.23298e-17
C3815	XI1/XI1/XI4/PHINOT#6	GND	2.42089e-17
C3816	XI1/XI0/XI0/ANOT#4	GND	9.81082e-18
C3817	XI1/XI0/XI0/ANOT#9	GND	4.88348e-17
C3818	XI1/XI0/XI0/ANOT#6	GND	1.02907e-17
C3819	VDD#31	GND	3.60805e-19
C3820	VDD#30	GND	1.26825e-18
C3821	XI1/XI1/D#6	GND	1.74398e-17
C3822	XI1/XI1/D#16	GND	2.45897e-17
C3823	VDD#165	GND	7.14874e-20
C3824	VDD#28	GND	8.37146e-19
C3825	VDD#126	GND	5.95395e-17
C3826	VDD#166	GND	4.90747e-17
C3827	net7#14	GND	2.8667e-17
C3828	net7#21	GND	8.96238e-17
C3829	SOUT0#18	GND	4.38955e-17
C3830	SOUT0#20	GND	6.30224e-17
C3831	SOUT0#22	GND	3.18348e-17
C3832	net7#12	GND	8.67498e-18
C3833	net7#15	GND	1.18863e-17
C3834	net7#10	GND	1.10923e-17
C3835	SOUT0#14	GND	3.23603e-18
C3836	SOUT0#19	GND	1.94159e-17
C3837	SOUT0#16	GND	8.43156e-18
C3838	VDD#26	GND	3.11409e-18
C3839	VDD#24	GND	2.60645e-19
C3840	VDD#170	GND	2.30328e-19
C3841	VDD#22	GND	2.25295e-18
C3842	XI0/net1#6	GND	3.57652e-19
C3843	XI0/XI0/XI0/BNOT#14	GND	9.80305e-18
C3844	XI0/XI0/XI0/BNOT#9	GND	3.07653e-17
C3845	XI0/XI0/XI0/BNOT#11	GND	1.8348e-17
C3846	XI0/XI0/XI1/net2#13	GND	1.75343e-17
C3847	XI0/XI0/XI1/net2#15	GND	2.92719e-17
C3848	XI0/net1#4	GND	6.20306e-18
C3849	XI0/net1#9	GND	7.68836e-18
C3850	XI0/net1#16	GND	2.01534e-17
C3851	XI0/XI1/XI4/net24#11	GND	2.17241e-18
C3852	XI0/XI1/XI4/net24#12	GND	1.17061e-17
C3853	XI0/XI1/Q#11	GND	2.17936e-17
C3854	XI0/XI1/Q#9	GND	1.09498e-17
C3855	XI0/XI0/XI1/net2#12	GND	8.07284e-18
C3856	VDD#20	GND	3.74949e-19
C3857	VDD#171	GND	3.8563e-19
C3858	VDD#18	GND	1.60408e-18
C3859	SOUT0#11	GND	1.47042e-17
C3860	SOUT0#24	GND	1.88875e-17
C3861	XI0/XI1/D#20	GND	3.08439e-18
C3862	XI0/XI1/D#17	GND	1.03658e-17
C3863	XI0/XI0/XI1/net2#16	GND	6.12784e-18
C3864	XI0/XI1/Q#6	GND	4.30485e-18
C3865	XI0/XI1/Q#12	GND	1.07738e-17
C3866	VDD#172	GND	2.20938e-19
C3867	VDD#16	GND	1.74327e-18
C3868	VDD#131	GND	2.81797e-20
C3869	VDD#14	GND	6.91838e-19
C3870	XI0/XI0/XI1/XI0/net13#4	GND	1.30885e-17
C3871	XI0/XI0/XI1/net2#9	GND	6.73319e-19
C3872	XI0/XI1/Q#5	GND	2.09121e-18
C3873	XI0/XI1/Q#7	GND	2.16707e-19
C3874	XI0/XI1/XI4/net24#13	GND	1.93822e-17
C3875	XI0/XI1/XI4/net24#6	GND	7.33241e-18
C3876	XI0/XI1/XI4/net24#9	GND	1.65682e-17
C3877	VDD#12	GND	6.90231e-19
C3878	XI0/XI1/D#19	GND	3.36909e-17
C3879	XI0/XI1/D#14	GND	2.50795e-17
C3880	CIN#11	GND	2.54602e-17
C3881	CIN#13	GND	4.17187e-17
C3882	VDD#10	GND	4.14886e-19
C3883	XI0/XI0/XI0/BNOT#5	GND	1.84278e-19
C3884	XI0/XI0/XI0/BNOT#10	GND	3.17641e-17
C3885	XI0/XI0/XI0/BNOT#7	GND	2.0708e-17
C3886	XI0/XI1/D#7	GND	8.64157e-19
C3887	XI0/XI1/XI5/net13#3	GND	1.06358e-17
C3888	VDD#175	GND	1.23331e-18
C3889	VDD#8	GND	2.68286e-19
C3890	XI0/XI1/D#15	GND	3.82381e-17
C3891	XI0/XI1/D#10	GND	6.97924e-18
C3892	XI0/XI1/XI4/PHINOT#4	GND	1.77609e-18
C3893	XI0/XI1/XI4/PHINOT#9	GND	5.23298e-17
C3894	XI0/XI1/XI4/PHINOT#6	GND	2.42089e-17
C3895	XI0/XI0/XI0/ANOT#4	GND	9.82796e-18
C3896	XI0/XI0/XI0/ANOT#9	GND	4.88217e-17
C3897	XI0/XI0/XI0/ANOT#6	GND	1.02907e-17
C3898	VDD#5	GND	3.60805e-19
C3899	VDD#4	GND	1.26825e-18
C3900	XI0/XI1/D#6	GND	1.74398e-17
C3901	XI0/XI1/D#16	GND	2.47453e-17
C3902	VDD#176	GND	7.14874e-20
C3903	VDD#2	GND	8.37146e-19
C3904	VDD#103	GND	3.24858e-19
C3905	VDD#85	GND	1.61383e-19
C3906	VDD#77	GND	3.24858e-19
C3907	VDD#59	GND	1.61383e-19
C3908	VDD#51	GND	3.24858e-19
C3909	VDD#33	GND	1.61383e-19
C3910	VDD#25	GND	3.24858e-19
C3911	VDD#7	GND	1.61383e-19
C3912	XI3/XI1/Q#8	GND	8.40992e-20
C3913	XI2/XI1/Q#8	GND	8.40992e-20
C3914	XI1/XI1/Q#8	GND	8.40992e-20
C3915	XI0/XI1/Q#8	GND	8.40992e-20
C3916	XI0/XI1/XI5/net13#5	GND	1.07128e-17
C3917	XI0/XI1/D#12	GND	5.19098e-18
C3918	XI0/XI0/XI1/XI0/net13#2	GND	1.40813e-17
C3919	XI0/XI0/XI1/net2#5	GND	1.61789e-18
C3920	XI0/net1#11	GND	3.5721e-19
C3921	XI0/net1#14	GND	8.13405e-18
C3922	XI0/net1#18	GND	6.35766e-18
C3923	XI1/XI1/XI5/net13#5	GND	1.07128e-17
C3924	XI1/XI1/D#12	GND	5.19098e-18
C3925	XI1/XI0/XI1/XI0/net13#2	GND	1.40813e-17
C3926	XI1/XI0/XI1/net2#5	GND	1.61789e-18
C3927	XI1/net1#11	GND	3.5721e-19
C3928	XI1/net1#14	GND	8.13405e-18
C3929	XI1/net1#18	GND	6.35766e-18
C3930	XI2/XI1/XI5/net13#5	GND	1.07128e-17
C3931	XI2/XI1/D#12	GND	5.19098e-18
C3932	XI2/XI0/XI1/XI0/net13#2	GND	1.40813e-17
C3933	XI2/XI0/XI1/net2#5	GND	1.61789e-18
C3934	XI2/net1#11	GND	3.5721e-19
C3935	XI2/net1#14	GND	8.13405e-18
C3936	XI2/net1#18	GND	6.35766e-18
C3937	XI3/XI1/XI5/net13#5	GND	1.07128e-17
C3938	XI3/XI1/D#12	GND	5.19098e-18
C3939	XI3/XI0/XI1/XI0/net13#2	GND	1.40813e-17
C3940	XI3/XI0/XI1/net2#5	GND	1.61789e-18
C3941	XI3/net1#11	GND	3.5721e-19
C3942	XI3/net1#14	GND	8.13405e-18
C3943	XI3/net1#18	GND	6.35766e-18
C3944	PHI#25	GND	5.02545e-17
C3945	RST#13	GND	9.43711e-17
*
*
.ENDS 4BIT_ACCUM
*
